//==============================================================================
//
// Project : MVP
//
// Verilog RTL(Behavioral) model
//
// This confidential and proprietary source code may be used only as authorized
// by a licensing agreement from ALPHAHOLDINGS Limited. The entire notice above
// must be reproduced on all authorized copies and copies may only be made to
// the extent permitted by a licensing agreement from ALPHAHOLDINGS Limited.
//
// COPYRIGHT (C) ALPHAHOLDINGS, inc. 2022
//
//==============================================================================
// File name : mvp1_hpdf
// Version : v1.1
// Description :
// Simulator : NC Verilog
// Created by : bhoh
// Date : 2023-12-14  16:18
//==============================================================================

module mvp1_hpdf (
    input              i_test_bypass,
    input              i_rstn_cpu2mvp,
    input              i_clk_cpu2mvp,
    input              i_clk_xtal_y,
    input              i_clk_mvp2main,
    input              i_clk_dvp4_y,
    input              i_clk_dvp5_y,
    input              i_clk_dvp6_y,
    input              i_clk_dvp7_y,
    input              i_clk_fcon,
    input              i_scan_clk,
    input              i_scan_mode,
    input              i_test_rstn,
    input   [  1:  0]  i_pll2551_mode,
    input   [  5:  0]  t_isp1_pll_p,
    input   [  9:  0]  t_isp1_pll_m,
    input   [  2:  0]  t_isp1_pll_s,
    input   [  1:  0]  t_isp1_pll_lock_con_in,
    input   [  1:  0]  t_isp1_pll_lock_con_out,
    input   [  1:  0]  t_isp1_pll_lock_con_dly,
    input   [  1:  0]  t_isp1_pll_lock_con_rev,
    input   [  4:  0]  t_isp1_pll_tst_afc,
    input   [  1:  0]  t_isp1_pll_icp,
    input              t_isp1_pll_resetb,
    input              t_isp1_pll_bypass,
    input              t_isp1_pll_tst_en,
    input              t_isp1_pll_fsel,
    input              t_isp1_pll_feed_en,
    input              t_isp1_pll_lock_en,
    input              t_isp1_pll_afcini_sel,
    input              t_isp1_pll_vcoini_en,
    input              t_isp1_pll_fout_mask,
    input              t_isp1_pll_pbias_ctrl,
    input              t_isp1_pll_pbias_ctrl_en,
    input   [  5:  0]  sr_isp1_pll_p,
    input   [  9:  0]  sr_isp1_pll_m,
    input   [  2:  0]  sr_isp1_pll_s,
    output             t_isp1_pll_feed_out,
    output             t_isp1_pll_lock,
    output             t_isp1_pll_fout,
    output             t_isp1_pll_sync_m_clk_out,
    output  [  4:  0]  t_isp1_pll_afc_code,
    output             o_irq_wdma_err_04,
    output             o_irq_wdma_err_05,
    output             o_irq_wdma_err_06,
    output             o_irq_wdma_err_07,
    output             o_irq_wdma_done_04,
    output             o_irq_wdma_done_05,
    output             o_irq_wdma_done_06,
    output             o_irq_wdma_done_07,
    output             o_irq_qisp1_0,
    output             o_irq_qisp1_1,
    input              i_isp4_cis_dvp_v_y,
    input              i_isp4_cis_dvp_h_y,
    input              i_isp4_cis_dvp_pv_y,
    input   [  9:  0]  i_isp4_cis_dvp_p_y,
    input              i_isp5_cis_dvp_v_y,
    input              i_isp5_cis_dvp_h_y,
    input              i_isp5_cis_dvp_pv_y,
    input   [  9:  0]  i_isp5_cis_dvp_p_y,
    input              i_isp6_cis_dvp_v_y,
    input              i_isp6_cis_dvp_h_y,
    input              i_isp6_cis_dvp_pv_y,
    input   [  9:  0]  i_isp6_cis_dvp_p_y,
    input              i_isp7_cis_dvp_v_y,
    input              i_isp7_cis_dvp_h_y,
    input              i_isp7_cis_dvp_pv_y,
    input   [  9:  0]  i_isp7_cis_dvp_p_y,
    input              i_test_mode,
    input   [ 38:  0]  i_ema,
    output             o_isp4_i2cm_scl_a,
    output             o_isp4_i2cm_scl_oe,
    input              i_isp4_i2cm_scl_y,
    output             o_isp4_i2cm_sda_a,
    output             o_isp4_i2cm_sda_oe,
    input              i_isp4_i2cm_sda_y,
    output             o_isp5_i2cm_scl_a,
    output             o_isp5_i2cm_scl_oe,
    input              i_isp5_i2cm_scl_y,
    output             o_isp5_i2cm_sda_a,
    output             o_isp5_i2cm_sda_oe,
    input              i_isp5_i2cm_sda_y,
    output             o_isp6_i2cm_scl_a,
    output             o_isp6_i2cm_scl_oe,
    input              i_isp6_i2cm_scl_y,
    output             o_isp6_i2cm_sda_a,
    output             o_isp6_i2cm_sda_oe,
    input              i_isp6_i2cm_sda_y,
    output             o_isp7_i2cm_scl_a,
    output             o_isp7_i2cm_scl_oe,
    input              i_isp7_i2cm_scl_y,
    output             o_isp7_i2cm_sda_a,
    output             o_isp7_i2cm_sda_oe,
    input              i_isp7_i2cm_sda_y,
    input              i_i2cs1_scl_y,
    output             o_i2cs1_sda_a,
    output             o_i2cs1_sda_oe,
    input              i_i2cs1_sda_y,
    input              i_mvp1_uart_rx_y,
    output             o_mvp1_uart_tx_a,
    output  [  9:  0]  o_isp4_cis_dvp_p_oe,
    output  [  9:  0]  o_isp5_cis_dvp_p_oe,
    output  [  9:  0]  o_isp6_cis_dvp_p_oe,
    output  [  9:  0]  o_isp7_cis_dvp_p_oe,
    output  [  9:  0]  o_isp4_cis_dvp_p_a,
    output  [  9:  0]  o_isp5_cis_dvp_p_a,
    output  [  9:  0]  o_isp6_cis_dvp_p_a,
    output  [  9:  0]  o_isp7_cis_dvp_p_a,
    output             o_isp4_cis_dvp_h_oe,
    output             o_isp5_cis_dvp_h_oe,
    output             o_isp6_cis_dvp_h_oe,
    output             o_isp7_cis_dvp_h_oe,
    output             o_isp4_cis_dvp_h_a,
    output             o_isp5_cis_dvp_h_a,
    output             o_isp6_cis_dvp_h_a,
    output             o_isp7_cis_dvp_h_a,
    output             o_isp4_cis_dvp_v_oe,
    output             o_isp5_cis_dvp_v_oe,
    output             o_isp6_cis_dvp_v_oe,
    output             o_isp7_cis_dvp_v_oe,
    output             o_isp4_cis_dvp_v_a,
    output             o_isp5_cis_dvp_v_a,
    output             o_isp6_cis_dvp_v_a,
    output             o_isp7_cis_dvp_v_a,
    input              MIPI_CLKP_RX4,
    input              MIPI_CLKN_RX4,
    input   [  3:  0]  MIPI_DP_RX4,
    input   [  3:  0]  MIPI_DN_RX4,
    input              MIPI_CLKP_RX5,
    input              MIPI_CLKN_RX5,
    input   [  3:  0]  MIPI_DP_RX5,
    input   [  3:  0]  MIPI_DN_RX5,
    input              MIPI_CLKP_RX6,
    input              MIPI_CLKN_RX6,
    input   [  3:  0]  MIPI_DP_RX6,
    input   [  3:  0]  MIPI_DN_RX6,
    input              MIPI_CLKP_RX7,
    input              MIPI_CLKN_RX7,
    input   [  3:  0]  MIPI_DP_RX7,
    input   [  3:  0]  MIPI_DN_RX7,
    input              MIPI_CHIP_EN_MR1,
    output             MIPI_HS_CKO_RX4,
    output  [  3:  0]  MIPI_HS_DO_RX4,
    output             MIPI_TEST_VMON_OUT_RX4,
    input              t_aclk,
    input              t_arstn,
    input              t_i2cs_scl,
    input              t_i_i2cs_sda,
    output             t_o_i2cs_sda,
    output             t_isp4_dvp_clk,
    output             t_isp4_dvp_v,
    output             t_isp4_dvp_h,
    output  [ 15:  0]  t_isp4_dvp_p,
    input              i_TM_7_MIPI_TEST,
    input   [  1:  0]  t_mipi_rx_test_sel,
    input              t_clk_isp4,
    input              t_clk_isp5,
    input              t_clk_isp6,
    input              t_clk_isp7,
    input              t_rstn_isp4,
    output             o_pix4_fstart,
    output             o_pix5_fstart,
    output             o_pix6_fstart,
    output             o_pix7_fstart,
    input              i_pix4_mask,
    input              i_pix5_mask,
    input              i_pix6_mask,
    input              i_pix7_mask,
    input              i_psel_cpu2mvp_1,
    input              i_penable_cpu2mvp_1,
    input              i_pwrite_cpu2mvp_1,
    input   [ 31:  0]  i_paddr_cpu2mvp_1,
    input   [ 31:  0]  i_pwdata_cpu2mvp_1,
    output             o_pready_cpu2mvp_1,
    output  [ 31:  0]  o_prdata_cpu2mvp_1,
    output             o_pslverr_cpu2mvp_1,
    output  [  1:  0]  o_awid_isp2main_1,
    output             o_awvalid_isp2main_1,
    input              i_awready_isp2main_1,
    output  [ 31:  0]  o_awaddr_isp2main_1,
    output  [  2:  0]  o_awprot_isp2main_1,
    output  [  7:  0]  o_awlen_isp2main_1,
    output  [  2:  0]  o_awsize_isp2main_1,
    output  [  1:  0]  o_awburst_isp2main_1,
    output             o_awlock_isp2main_1,
    output  [  3:  0]  o_awcache_isp2main_1,
    output             o_wvalid_isp2main_1,
    input              i_wready_isp2main_1,
    output  [127:  0]  o_wdata_isp2main_1,
    output  [ 15:  0]  o_wstrb_isp2main_1,
    output             o_wlast_isp2main_1,
    input   [  1:  0]  i_bid_isp2main_1,
    input              i_bvalid_isp2main_1,
    output             o_bready_isp2main_1,
    input   [  1:  0]  i_bresp_isp2main_1,
    output  [  1:  0]  o_arid_isp2main_1,
    output  [  2:  0]  o_arprot_isp2main_1,
    output             o_arvalid_isp2main_1,
    input              i_arready_isp2main_1,
    output  [ 31:  0]  o_araddr_isp2main_1,
    output  [  7:  0]  o_arlen_isp2main_1,
    output  [  2:  0]  o_arsize_isp2main_1,
    output  [  1:  0]  o_arburst_isp2main_1,
    output             o_arlock_isp2main_1,
    output  [  3:  0]  o_arcache_isp2main_1,
    input   [  1:  0]  i_rid_isp2main_1,
    input              i_rvalid_isp2main_1,
    output             o_rready_isp2main_1,
    input   [127:  0]  i_rdata_isp2main_1,
    input              i_rlast_isp2main_1,
    input   [  1:  0]  i_rresp_isp2main_1,
    output  [  1:  0]  o_awuser_isp2main_1,
    output  [  1:  0]  o_aruser_isp2main_1
);

    wire            mvp1_crm_o_pll_isp1_norm_resetb;
    wire            mvp1_crm_o_pll_isp1_norm_bypass;
    wire    [ 5:0]  mvp1_crm_o_pll_isp1_norm_p;
    wire    [ 9:0]  mvp1_crm_o_pll_isp1_norm_m;
    wire    [ 2:0]  mvp1_crm_o_pll_isp1_norm_s;
    wire            mvp1_crm_o_pll_isp1_norm_lock_en;
    wire    [ 1:0]  mvp1_crm_o_pll_isp1_norm_lock_con_in;
    wire    [ 1:0]  mvp1_crm_o_pll_isp1_norm_lock_con_out;
    wire    [ 1:0]  mvp1_crm_o_pll_isp1_norm_lock_con_dly;
    wire    [ 1:0]  mvp1_crm_o_pll_isp1_norm_lock_con_rev;
    wire            mvp1_crm_o_pll_isp1_norm_feed_en;
    wire            mvp1_crm_o_pll_isp1_norm_fsel;
    wire            mvp1_crm_o_pll_isp1_norm_tst_en;
    wire    [ 4:0]  mvp1_crm_o_pll_isp1_norm_tst_afc;
    wire            mvp1_crm_o_pll_isp1_norm_afcini_sel;
    wire            mvp1_crm_o_pll_isp1_norm_vcoini_en;
    wire            mvp1_crm_o_pll_isp1_norm_fout_mask;
    wire            mvp1_crm_o_pll_isp1_norm_pbias_ctrl;
    wire            mvp1_crm_o_pll_isp1_norm_pbias_ctrl_en;
    wire    [ 1:0]  mvp1_crm_o_pll_isp1_norm_icp;
    wire            mvp1_crm_o_clk_phy_ref;
    wire            mvp1_crm_o_clk_riscv_timer1;
    wire            mvp1_crm_o_rstn_riscv_timer1;
    wire            mvp1_crm_o_clk_cpu2mvp;
    wire            mvp1_crm_o_rstn_cpu2mvp;
    wire            mvp1_crm_o_sclk_wdma4;
    wire            mvp1_crm_o_srstn_wdma4;
    wire            mvp1_crm_o_sclk_wdma5;
    wire            mvp1_crm_o_srstn_wdma5;
    wire            mvp1_crm_o_sclk_wdma6;
    wire            mvp1_crm_o_srstn_wdma6;
    wire            mvp1_crm_o_sclk_wdma7;
    wire            mvp1_crm_o_srstn_wdma7;
    wire            mvp1_crm_o_clk_fcon1;
    wire            mvp1_crm_o_rstn_fcon1;
    wire            mvp1_crm_o_clk_mvp2main;
    wire            mvp1_crm_o_rstn_mvp2main;
    wire            mvp1_crm_o_mclk_wdma4;
    wire            mvp1_crm_o_mrstn_wdma4;
    wire            mvp1_crm_o_mclk_wdma5;
    wire            mvp1_crm_o_mrstn_wdma5;
    wire            mvp1_crm_o_mclk_wdma6;
    wire            mvp1_crm_o_mrstn_wdma6;
    wire            mvp1_crm_o_mclk_wdma7;
    wire            mvp1_crm_o_mrstn_wdma7;
    wire            mvp1_crm_o_clk_riscv;
    wire            mvp1_crm_o_rstn_riscv;
    wire            mvp1_crm_o_clk_dvp4;
    wire            mvp1_crm_o_rstn_dvp4;
    wire            mvp1_crm_o_clk_dvp5;
    wire            mvp1_crm_o_rstn_dvp5;
    wire            mvp1_crm_o_clk_dvp6;
    wire            mvp1_crm_o_rstn_dvp6;
    wire            mvp1_crm_o_clk_dvp7;
    wire            mvp1_crm_o_rstn_dvp7;
    wire            mvp1_crm_o_clk_isp4_clk;
    wire            mvp1_crm_o_rstn_isp4_clk;
    wire            mvp1_crm_o_clk_isp5_clk;
    wire            mvp1_crm_o_rstn_isp5_clk;
    wire            mvp1_crm_o_clk_isp6_clk;
    wire            mvp1_crm_o_rstn_isp6_clk;
    wire            mvp1_crm_o_clk_isp7_clk;
    wire            mvp1_crm_o_rstn_isp7_clk;
    wire            mvp1_crm_o_rstn_isp4;
    wire            mvp1_crm_o_rstn_isp5;
    wire            mvp1_crm_o_rstn_isp6;
    wire            mvp1_crm_o_rstn_isp7;
    wire            isp1_pll_o_feed_out;
    wire            isp1_pll_o_lock;
    wire            isp1_pll_o_fout;
    wire            isp1_pll_o_sync_m_clk_out;
    wire    [ 4:0]  isp1_pll_o_afc_code;
    wire            mvp1_sub_o_isp4_clk;
    wire            mvp1_sub_o_isp5_clk;
    wire            mvp1_sub_o_isp6_clk;
    wire            mvp1_sub_o_isp7_clk;
    wire            mvp1_sub_o_mvp1_crm_psel;
    wire            mvp1_sub_o_mvp1_crm_penable;
    wire            mvp1_sub_o_mvp1_crm_pwrite;
    wire    [11:0]  mvp1_sub_o_mvp1_crm_paddr;
    wire    [31:0]  mvp1_sub_o_mvp1_crm_pwdata;
    wire    [31:0]  mvp1_sub_i_mvp1_crm_prdata;

    assign  t_isp1_pll_afc_code[4:0] = isp1_pll_o_afc_code[4:0];
    assign  t_isp1_pll_feed_out = isp1_pll_o_feed_out;
    assign  t_isp1_pll_fout = isp1_pll_o_fout;
    assign  t_isp1_pll_lock = isp1_pll_o_lock;
    assign  t_isp1_pll_sync_m_clk_out = isp1_pll_o_sync_m_clk_out;

    mvp_crm_mvp1 u_mvp1_crm (
        .i_test_bypass                   (i_test_bypass),
        .i_rstn_mvp                      (i_rstn_cpu2mvp),
        .i_apb_pclk                      (i_clk_cpu2mvp),
        .i_apb_prstn                     (i_rstn_cpu2mvp),
        .i_apb_psel                      (mvp1_sub_o_mvp1_crm_psel),
        .i_apb_penable                   (mvp1_sub_o_mvp1_crm_penable),
        .i_apb_pwrite                    (mvp1_sub_o_mvp1_crm_pwrite),
        .i_apb_paddr                     (mvp1_sub_o_mvp1_crm_paddr),
        .i_apb_pwdata                    (mvp1_sub_o_mvp1_crm_pwdata),
        .o_apb_prdata                    (mvp1_sub_i_mvp1_crm_prdata),
        .o_pll_isp1_norm_resetb          (mvp1_crm_o_pll_isp1_norm_resetb),
        .o_pll_isp1_norm_bypass          (mvp1_crm_o_pll_isp1_norm_bypass),
        .o_pll_isp1_norm_p               (mvp1_crm_o_pll_isp1_norm_p),
        .o_pll_isp1_norm_m               (mvp1_crm_o_pll_isp1_norm_m),
        .o_pll_isp1_norm_s               (mvp1_crm_o_pll_isp1_norm_s),
        .i_pll_isp1_lock                 (isp1_pll_o_lock),
        .i_pll_isp1_feed_out             (isp1_pll_o_feed_out),
        .i_pll_isp1_sync_m_clk_out       (isp1_pll_o_sync_m_clk_out),
        .i_pll_isp1_afc_code             (isp1_pll_o_afc_code),
        .o_pll_isp1_norm_lock_en         (mvp1_crm_o_pll_isp1_norm_lock_en),
        .o_pll_isp1_norm_lock_con_in     (mvp1_crm_o_pll_isp1_norm_lock_con_in),
        .o_pll_isp1_norm_lock_con_out    (mvp1_crm_o_pll_isp1_norm_lock_con_out),
        .o_pll_isp1_norm_lock_con_dly    (mvp1_crm_o_pll_isp1_norm_lock_con_dly),
        .o_pll_isp1_norm_lock_con_rev    (mvp1_crm_o_pll_isp1_norm_lock_con_rev),
        .o_pll_isp1_norm_feed_en         (mvp1_crm_o_pll_isp1_norm_feed_en),
        .o_pll_isp1_norm_fsel            (mvp1_crm_o_pll_isp1_norm_fsel),
        .o_pll_isp1_norm_tst_en          (mvp1_crm_o_pll_isp1_norm_tst_en),
        .o_pll_isp1_norm_tst_afc         (mvp1_crm_o_pll_isp1_norm_tst_afc),
        .o_pll_isp1_norm_afcini_sel      (mvp1_crm_o_pll_isp1_norm_afcini_sel),
        .o_pll_isp1_norm_vcoini_en       (mvp1_crm_o_pll_isp1_norm_vcoini_en),
        .o_pll_isp1_norm_fout_mask       (mvp1_crm_o_pll_isp1_norm_fout_mask),
        .o_pll_isp1_norm_pbias_ctrl      (mvp1_crm_o_pll_isp1_norm_pbias_ctrl),
        .o_pll_isp1_norm_pbias_ctrl_en   (mvp1_crm_o_pll_isp1_norm_pbias_ctrl_en),
        .o_pll_isp1_norm_icp             (mvp1_crm_o_pll_isp1_norm_icp),
        .i_clk_xtal_y                    (i_clk_xtal_y),
        .i_clk_cpu2mvp                   (i_clk_cpu2mvp),
        .i_clk_mvp2main                  (i_clk_mvp2main),
        .i_clk_dvp4_y                    (i_clk_dvp4_y),
        .i_clk_dvp5_y                    (i_clk_dvp5_y),
        .i_clk_dvp6_y                    (i_clk_dvp6_y),
        .i_clk_dvp7_y                    (i_clk_dvp7_y),
        .i_pll_isp1                      (isp1_pll_o_fout),
        .i_clk_fcon                      (i_clk_fcon),
        .i_clk_isp4                      (mvp1_sub_o_isp4_clk),
        .i_clk_isp5                      (mvp1_sub_o_isp5_clk),
        .i_clk_isp6                      (mvp1_sub_o_isp6_clk),
        .i_clk_isp7                      (mvp1_sub_o_isp7_clk),
        .o_clk_phy_ref                   (mvp1_crm_o_clk_phy_ref),
        .o_clk_riscv_timer1              (mvp1_crm_o_clk_riscv_timer1),
        .o_rstn_riscv_timer1             (mvp1_crm_o_rstn_riscv_timer1),
        .o_clk_cpu2mvp                   (mvp1_crm_o_clk_cpu2mvp),
        .o_rstn_cpu2mvp                  (mvp1_crm_o_rstn_cpu2mvp),
        .o_sclk_wdma4                    (mvp1_crm_o_sclk_wdma4),
        .o_srstn_wdma4                   (mvp1_crm_o_srstn_wdma4),
        .o_sclk_wdma5                    (mvp1_crm_o_sclk_wdma5),
        .o_srstn_wdma5                   (mvp1_crm_o_srstn_wdma5),
        .o_sclk_wdma6                    (mvp1_crm_o_sclk_wdma6),
        .o_srstn_wdma6                   (mvp1_crm_o_srstn_wdma6),
        .o_sclk_wdma7                    (mvp1_crm_o_sclk_wdma7),
        .o_srstn_wdma7                   (mvp1_crm_o_srstn_wdma7),
        .o_clk_fcon1                     (mvp1_crm_o_clk_fcon1),
        .o_rstn_fcon1                    (mvp1_crm_o_rstn_fcon1),
        .o_clk_mvp2main                  (mvp1_crm_o_clk_mvp2main),
        .o_rstn_mvp2main                 (mvp1_crm_o_rstn_mvp2main),
        .o_mclk_wdma4                    (mvp1_crm_o_mclk_wdma4),
        .o_mrstn_wdma4                   (mvp1_crm_o_mrstn_wdma4),
        .o_mclk_wdma5                    (mvp1_crm_o_mclk_wdma5),
        .o_mrstn_wdma5                   (mvp1_crm_o_mrstn_wdma5),
        .o_mclk_wdma6                    (mvp1_crm_o_mclk_wdma6),
        .o_mrstn_wdma6                   (mvp1_crm_o_mrstn_wdma6),
        .o_mclk_wdma7                    (mvp1_crm_o_mclk_wdma7),
        .o_mrstn_wdma7                   (mvp1_crm_o_mrstn_wdma7),
        .o_clk_riscv                     (mvp1_crm_o_clk_riscv),
        .o_rstn_riscv                    (mvp1_crm_o_rstn_riscv),
        .o_clk_dvp4                      (mvp1_crm_o_clk_dvp4),
        .o_rstn_dvp4                     (mvp1_crm_o_rstn_dvp4),
        .o_clk_dvp5                      (mvp1_crm_o_clk_dvp5),
        .o_rstn_dvp5                     (mvp1_crm_o_rstn_dvp5),
        .o_clk_dvp6                      (mvp1_crm_o_clk_dvp6),
        .o_rstn_dvp6                     (mvp1_crm_o_rstn_dvp6),
        .o_clk_dvp7                      (mvp1_crm_o_clk_dvp7),
        .o_rstn_dvp7                     (mvp1_crm_o_rstn_dvp7),
        .o_clk_isp4_clk                  (mvp1_crm_o_clk_isp4_clk),
        .o_rstn_isp4_clk                 (mvp1_crm_o_rstn_isp4_clk),
        .o_clk_isp5_clk                  (mvp1_crm_o_clk_isp5_clk),
        .o_rstn_isp5_clk                 (mvp1_crm_o_rstn_isp5_clk),
        .o_clk_isp6_clk                  (mvp1_crm_o_clk_isp6_clk),
        .o_rstn_isp6_clk                 (mvp1_crm_o_rstn_isp6_clk),
        .o_clk_isp7_clk                  (mvp1_crm_o_clk_isp7_clk),
        .o_rstn_isp7_clk                 (mvp1_crm_o_rstn_isp7_clk),
        .o_rstn_isp4                     (mvp1_crm_o_rstn_isp4),
        .o_rstn_isp5                     (mvp1_crm_o_rstn_isp5),
        .o_rstn_isp6                     (mvp1_crm_o_rstn_isp6),
        .o_rstn_isp7                     (mvp1_crm_o_rstn_isp7),
        .i_scan_clk                      (i_scan_clk),
        .i_scan_mode                     (i_scan_mode),
        .i_scan_rstn                     (i_test_rstn)
    );

    tmux_sf_pll2551x_ln28lpp_5000 u_pll_isp1 (
        .i_tmode                         (i_pll2551_mode),
        .i_norm_p                        (mvp1_crm_o_pll_isp1_norm_p),
        .i_norm_m                        (mvp1_crm_o_pll_isp1_norm_m),
        .i_norm_s                        (mvp1_crm_o_pll_isp1_norm_s),
        .i_norm_lock_con_in              (mvp1_crm_o_pll_isp1_norm_lock_con_in),
        .i_norm_lock_con_out             (mvp1_crm_o_pll_isp1_norm_lock_con_out),
        .i_norm_lock_con_dly             (mvp1_crm_o_pll_isp1_norm_lock_con_dly),
        .i_norm_lock_con_rev             (mvp1_crm_o_pll_isp1_norm_lock_con_rev),
        .i_norm_tst_afc                  (mvp1_crm_o_pll_isp1_norm_tst_afc),
        .i_norm_icp                      (mvp1_crm_o_pll_isp1_norm_icp),
        .i_norm_fin                      (mvp1_crm_o_clk_phy_ref),
        .i_norm_resetb                   (mvp1_crm_o_pll_isp1_norm_resetb),
        .i_norm_bypass                   (mvp1_crm_o_pll_isp1_norm_bypass),
        .i_norm_tst_en                   (mvp1_crm_o_pll_isp1_norm_tst_en),
        .i_norm_fsel                     (mvp1_crm_o_pll_isp1_norm_fsel),
        .i_norm_feed_en                  (mvp1_crm_o_pll_isp1_norm_feed_en),
        .i_norm_lock_en                  (mvp1_crm_o_pll_isp1_norm_lock_en),
        .i_norm_afcini_sel               (mvp1_crm_o_pll_isp1_norm_afcini_sel),
        .i_norm_vcoini_en                (mvp1_crm_o_pll_isp1_norm_vcoini_en),
        .i_norm_fout_mask                (mvp1_crm_o_pll_isp1_norm_fout_mask),
        .i_norm_pbias_ctrl               (mvp1_crm_o_pll_isp1_norm_pbias_ctrl),
        .i_norm_pbias_ctrl_en            (mvp1_crm_o_pll_isp1_norm_pbias_ctrl_en),
        .i_test0_p                       (t_isp1_pll_p),
        .i_test0_m                       (t_isp1_pll_m),
        .i_test0_s                       (t_isp1_pll_s),
        .i_test0_lock_con_in             (t_isp1_pll_lock_con_in),
        .i_test0_lock_con_out            (t_isp1_pll_lock_con_out),
        .i_test0_lock_con_dly            (t_isp1_pll_lock_con_dly),
        .i_test0_lock_con_rev            (t_isp1_pll_lock_con_rev),
        .i_test0_tst_afc                 (t_isp1_pll_tst_afc),
        .i_test0_icp                     (t_isp1_pll_icp),
        .i_test0_fin                     (i_clk_xtal_y),
        .i_test0_resetb                  (t_isp1_pll_resetb),
        .i_test0_bypass                  (t_isp1_pll_bypass),
        .i_test0_tst_en                  (t_isp1_pll_tst_en),
        .i_test0_fsel                    (t_isp1_pll_fsel),
        .i_test0_feed_en                 (t_isp1_pll_feed_en),
        .i_test0_lock_en                 (t_isp1_pll_lock_en),
        .i_test0_afcini_sel              (t_isp1_pll_afcini_sel),
        .i_test0_vcoini_en               (t_isp1_pll_vcoini_en),
        .i_test0_fout_mask               (t_isp1_pll_fout_mask),
        .i_test0_pbias_ctrl              (t_isp1_pll_pbias_ctrl),
        .i_test0_pbias_ctrl_en           (t_isp1_pll_pbias_ctrl_en),
        .i_test1_p                       (sr_isp1_pll_p),
        .i_test1_m                       (sr_isp1_pll_m),
        .i_test1_s                       (sr_isp1_pll_s),
        .i_test1_lock_con_in             (2'h3),
        .i_test1_lock_con_out            (2'h3),
        .i_test1_lock_con_dly            (2'h3),
        .i_test1_lock_con_rev            (2'h0),
        .i_test1_tst_afc                 (5'h0),
        .i_test1_icp                     (2'h0),
        .i_test1_fin                     (i_clk_xtal_y),
        .i_test1_resetb                  (t_isp1_pll_resetb),
        .i_test1_bypass                  (1'h0),
        .i_test1_tst_en                  (1'h0),
        .i_test1_fsel                    (1'h0),
        .i_test1_feed_en                 (1'h0),
        .i_test1_lock_en                 (1'h1),
        .i_test1_afcini_sel              (1'h0),
        .i_test1_vcoini_en               (1'h1),
        .i_test1_fout_mask               (1'h0),
        .i_test1_pbias_ctrl              (1'h0),
        .i_test1_pbias_ctrl_en           (1'h0),
        .o_feed_out                      (isp1_pll_o_feed_out),
        .o_lock                          (isp1_pll_o_lock),
        .o_fout                          (isp1_pll_o_fout),
        .o_sync_m_clk_out                (isp1_pll_o_sync_m_clk_out),
        .o_afc_code                      (isp1_pll_o_afc_code)
    );

    mvp1_sub u_mvp1_sub (
        .i_clk_phy_ref                   (mvp1_crm_o_clk_phy_ref),
        .i_clk_riscv_timer1              (mvp1_crm_o_clk_riscv_timer1),
        .i_rstn_riscv_timer1             (mvp1_crm_o_rstn_riscv_timer1),
        .i_clk_cpu2mvp                   (mvp1_crm_o_clk_cpu2mvp),
        .i_rstn_cpu2mvp                  (mvp1_crm_o_rstn_cpu2mvp),
        .i_sclk_wdma4                    (mvp1_crm_o_sclk_wdma4),
        .i_srstn_wdma4                   (mvp1_crm_o_srstn_wdma4),
        .i_sclk_wdma5                    (mvp1_crm_o_sclk_wdma5),
        .i_srstn_wdma5                   (mvp1_crm_o_srstn_wdma5),
        .i_sclk_wdma6                    (mvp1_crm_o_sclk_wdma6),
        .i_srstn_wdma6                   (mvp1_crm_o_srstn_wdma6),
        .i_sclk_wdma7                    (mvp1_crm_o_sclk_wdma7),
        .i_srstn_wdma7                   (mvp1_crm_o_srstn_wdma7),
        .i_clk_mvp2main                  (mvp1_crm_o_clk_mvp2main),
        .i_rstn_mvp2main                 (mvp1_crm_o_rstn_mvp2main),
        .i_mclk_wdma4                    (mvp1_crm_o_mclk_wdma4),
        .i_mrstn_wdma4                   (mvp1_crm_o_mrstn_wdma4),
        .i_mclk_wdma5                    (mvp1_crm_o_mclk_wdma5),
        .i_mrstn_wdma5                   (mvp1_crm_o_mrstn_wdma5),
        .i_mclk_wdma6                    (mvp1_crm_o_mclk_wdma6),
        .i_mrstn_wdma6                   (mvp1_crm_o_mrstn_wdma6),
        .i_mclk_wdma7                    (mvp1_crm_o_mclk_wdma7),
        .i_mrstn_wdma7                   (mvp1_crm_o_mrstn_wdma7),
        .i_clk_riscv                     (mvp1_crm_o_clk_riscv),
        .i_rstn_riscv                    (mvp1_crm_o_rstn_riscv),
        .i_clk_dvp4_y                    (mvp1_crm_o_clk_dvp4),
        .i_rstn_dvp4_y                   (mvp1_crm_o_rstn_dvp4),
        .i_clk_dvp5_y                    (mvp1_crm_o_clk_dvp5),
        .i_rstn_dvp5_y                   (mvp1_crm_o_rstn_dvp5),
        .i_clk_dvp6_y                    (mvp1_crm_o_clk_dvp6),
        .i_rstn_dvp6_y                   (mvp1_crm_o_rstn_dvp6),
        .i_clk_dvp7_y                    (mvp1_crm_o_clk_dvp7),
        .i_rstn_dvp7_y                   (mvp1_crm_o_rstn_dvp7),
        .i_clk_isp4                      (mvp1_crm_o_clk_isp4_clk),
        .i_rstn_isp4                     (mvp1_crm_o_rstn_isp4_clk),
        .i_clk_isp5                      (mvp1_crm_o_clk_isp5_clk),
        .i_rstn_isp5                     (mvp1_crm_o_rstn_isp5_clk),
        .i_clk_isp6                      (mvp1_crm_o_clk_isp6_clk),
        .i_rstn_isp6                     (mvp1_crm_o_rstn_isp6_clk),
        .i_clk_isp7                      (mvp1_crm_o_clk_isp7_clk),
        .i_rstn_isp7                     (mvp1_crm_o_rstn_isp7_clk),
        .i_clk_fcon1                     (mvp1_crm_o_clk_fcon1),
        .i_rstn_fcon1                    (mvp1_crm_o_rstn_fcon1),
        .o_isp4_clk                      (mvp1_sub_o_isp4_clk),
        .o_isp5_clk                      (mvp1_sub_o_isp5_clk),
        .o_isp6_clk                      (mvp1_sub_o_isp6_clk),
        .o_isp7_clk                      (mvp1_sub_o_isp7_clk),
        .i_isp4_rstn                     (mvp1_crm_o_rstn_isp4),
        .i_isp5_rstn                     (mvp1_crm_o_rstn_isp5),
        .i_isp6_rstn                     (mvp1_crm_o_rstn_isp6),
        .i_isp7_rstn                     (mvp1_crm_o_rstn_isp7),
        .o_irq_wdma_err_04               (o_irq_wdma_err_04),
        .o_irq_wdma_err_05               (o_irq_wdma_err_05),
        .o_irq_wdma_err_06               (o_irq_wdma_err_06),
        .o_irq_wdma_err_07               (o_irq_wdma_err_07),
        .o_irq_wdma_done_04              (o_irq_wdma_done_04),
        .o_irq_wdma_done_05              (o_irq_wdma_done_05),
        .o_irq_wdma_done_06              (o_irq_wdma_done_06),
        .o_irq_wdma_done_07              (o_irq_wdma_done_07),
        .o_irq_qisp1_0                   (o_irq_qisp1_0),
        .o_irq_qisp1_1                   (o_irq_qisp1_1),
        .i_psel_cpu2mvp_1                (i_psel_cpu2mvp_1),
        .i_penable_cpu2mvp_1             (i_penable_cpu2mvp_1),
        .i_pwrite_cpu2mvp_1              (i_pwrite_cpu2mvp_1),
        .i_paddr_cpu2mvp_1               (i_paddr_cpu2mvp_1),
        .i_pwdata_cpu2mvp_1              (i_pwdata_cpu2mvp_1),
        .o_pready_cpu2mvp_1              (o_pready_cpu2mvp_1),
        .o_prdata_cpu2mvp_1              (o_prdata_cpu2mvp_1),
        .o_pslverr_cpu2mvp_1             (o_pslverr_cpu2mvp_1),
        .o_awid_isp2main_1               (o_awid_isp2main_1),
        .o_awvalid_isp2main_1            (o_awvalid_isp2main_1),
        .i_awready_isp2main_1            (i_awready_isp2main_1),
        .o_awaddr_isp2main_1             (o_awaddr_isp2main_1),
        .o_awprot_isp2main_1             (o_awprot_isp2main_1),
        .o_awlen_isp2main_1              (o_awlen_isp2main_1),
        .o_awsize_isp2main_1             (o_awsize_isp2main_1),
        .o_awburst_isp2main_1            (o_awburst_isp2main_1),
        .o_awlock_isp2main_1             (o_awlock_isp2main_1),
        .o_awcache_isp2main_1            (o_awcache_isp2main_1),
        .o_wvalid_isp2main_1             (o_wvalid_isp2main_1),
        .i_wready_isp2main_1             (i_wready_isp2main_1),
        .o_wdata_isp2main_1              (o_wdata_isp2main_1),
        .o_wstrb_isp2main_1              (o_wstrb_isp2main_1),
        .o_wlast_isp2main_1              (o_wlast_isp2main_1),
        .i_bid_isp2main_1                (i_bid_isp2main_1),
        .i_bvalid_isp2main_1             (i_bvalid_isp2main_1),
        .o_bready_isp2main_1             (o_bready_isp2main_1),
        .i_bresp_isp2main_1              (i_bresp_isp2main_1),
        .o_arid_isp2main_1               (o_arid_isp2main_1),
        .o_arprot_isp2main_1             (o_arprot_isp2main_1),
        .o_arvalid_isp2main_1            (o_arvalid_isp2main_1),
        .i_arready_isp2main_1            (i_arready_isp2main_1),
        .o_araddr_isp2main_1             (o_araddr_isp2main_1),
        .o_arlen_isp2main_1              (o_arlen_isp2main_1),
        .o_arsize_isp2main_1             (o_arsize_isp2main_1),
        .o_arburst_isp2main_1            (o_arburst_isp2main_1),
        .o_arlock_isp2main_1             (o_arlock_isp2main_1),
        .o_arcache_isp2main_1            (o_arcache_isp2main_1),
        .i_rid_isp2main_1                (i_rid_isp2main_1),
        .i_rvalid_isp2main_1             (i_rvalid_isp2main_1),
        .o_rready_isp2main_1             (o_rready_isp2main_1),
        .i_rdata_isp2main_1              (i_rdata_isp2main_1),
        .i_rlast_isp2main_1              (i_rlast_isp2main_1),
        .i_rresp_isp2main_1              (i_rresp_isp2main_1),
        .o_mvp1_crm_psel                 (mvp1_sub_o_mvp1_crm_psel),
        .o_mvp1_crm_penable              (mvp1_sub_o_mvp1_crm_penable),
        .o_mvp1_crm_pwrite               (mvp1_sub_o_mvp1_crm_pwrite),
        .o_mvp1_crm_paddr                (mvp1_sub_o_mvp1_crm_paddr),
        .o_mvp1_crm_pwdata               (mvp1_sub_o_mvp1_crm_pwdata),
        .i_mvp1_crm_prdata               (mvp1_sub_i_mvp1_crm_prdata),
        .i_mvp1_crm_pready               (1'h1),
        .i_mvp1_crm_pslverr              (1'h0),
        .i_isp4_cis_dvp_v_y              (i_isp4_cis_dvp_v_y),
        .i_isp4_cis_dvp_h_y              (i_isp4_cis_dvp_h_y),
        .i_isp4_cis_dvp_pv_y             (i_isp4_cis_dvp_pv_y),
        .i_isp4_cis_dvp_p_y              (i_isp4_cis_dvp_p_y),
        .i_isp5_cis_dvp_v_y              (i_isp5_cis_dvp_v_y),
        .i_isp5_cis_dvp_h_y              (i_isp5_cis_dvp_h_y),
        .i_isp5_cis_dvp_pv_y             (i_isp5_cis_dvp_pv_y),
        .i_isp5_cis_dvp_p_y              (i_isp5_cis_dvp_p_y),
        .i_isp6_cis_dvp_v_y              (i_isp6_cis_dvp_v_y),
        .i_isp6_cis_dvp_h_y              (i_isp6_cis_dvp_h_y),
        .i_isp6_cis_dvp_pv_y             (i_isp6_cis_dvp_pv_y),
        .i_isp6_cis_dvp_p_y              (i_isp6_cis_dvp_p_y),
        .i_isp7_cis_dvp_v_y              (i_isp7_cis_dvp_v_y),
        .i_isp7_cis_dvp_h_y              (i_isp7_cis_dvp_h_y),
        .i_isp7_cis_dvp_pv_y             (i_isp7_cis_dvp_pv_y),
        .i_isp7_cis_dvp_p_y              (i_isp7_cis_dvp_p_y),
        .i_test_mode                     (i_test_mode),
        .i_test_bypass                   (i_test_bypass),
        .i_ema                           (i_ema),
        .o_isp4_i2cm_scl_a               (o_isp4_i2cm_scl_a),
        .o_isp4_i2cm_scl_oe              (o_isp4_i2cm_scl_oe),
        .i_isp4_i2cm_scl_y               (i_isp4_i2cm_scl_y),
        .o_isp4_i2cm_sda_a               (o_isp4_i2cm_sda_a),
        .o_isp4_i2cm_sda_oe              (o_isp4_i2cm_sda_oe),
        .i_isp4_i2cm_sda_y               (i_isp4_i2cm_sda_y),
        .o_isp5_i2cm_scl_a               (o_isp5_i2cm_scl_a),
        .o_isp5_i2cm_scl_oe              (o_isp5_i2cm_scl_oe),
        .i_isp5_i2cm_scl_y               (i_isp5_i2cm_scl_y),
        .o_isp5_i2cm_sda_a               (o_isp5_i2cm_sda_a),
        .o_isp5_i2cm_sda_oe              (o_isp5_i2cm_sda_oe),
        .i_isp5_i2cm_sda_y               (i_isp5_i2cm_sda_y),
        .o_isp6_i2cm_scl_a               (o_isp6_i2cm_scl_a),
        .o_isp6_i2cm_scl_oe              (o_isp6_i2cm_scl_oe),
        .i_isp6_i2cm_scl_y               (i_isp6_i2cm_scl_y),
        .o_isp6_i2cm_sda_a               (o_isp6_i2cm_sda_a),
        .o_isp6_i2cm_sda_oe              (o_isp6_i2cm_sda_oe),
        .i_isp6_i2cm_sda_y               (i_isp6_i2cm_sda_y),
        .o_isp7_i2cm_scl_a               (o_isp7_i2cm_scl_a),
        .o_isp7_i2cm_scl_oe              (o_isp7_i2cm_scl_oe),
        .i_isp7_i2cm_scl_y               (i_isp7_i2cm_scl_y),
        .o_isp7_i2cm_sda_a               (o_isp7_i2cm_sda_a),
        .o_isp7_i2cm_sda_oe              (o_isp7_i2cm_sda_oe),
        .i_isp7_i2cm_sda_y               (i_isp7_i2cm_sda_y),
        .i_i2cs1_scl_y                   (i_i2cs1_scl_y),
        .o_i2cs1_sda_a                   (o_i2cs1_sda_a),
        .o_i2cs1_sda_oe                  (o_i2cs1_sda_oe),
        .i_i2cs1_sda_y                   (i_i2cs1_sda_y),
        .i_mvp1_uart_rx_y                (i_mvp1_uart_rx_y),
        .o_mvp1_uart_tx_a                (o_mvp1_uart_tx_a),
        .o_isp4_cis_dvp_p_oe             (o_isp4_cis_dvp_p_oe),
        .o_isp5_cis_dvp_p_oe             (o_isp5_cis_dvp_p_oe),
        .o_isp6_cis_dvp_p_oe             (o_isp6_cis_dvp_p_oe),
        .o_isp7_cis_dvp_p_oe             (o_isp7_cis_dvp_p_oe),
        .o_isp4_cis_dvp_p_a              (o_isp4_cis_dvp_p_a),
        .o_isp5_cis_dvp_p_a              (o_isp5_cis_dvp_p_a),
        .o_isp6_cis_dvp_p_a              (o_isp6_cis_dvp_p_a),
        .o_isp7_cis_dvp_p_a              (o_isp7_cis_dvp_p_a),
        .o_isp4_cis_dvp_h_oe             (o_isp4_cis_dvp_h_oe),
        .o_isp5_cis_dvp_h_oe             (o_isp5_cis_dvp_h_oe),
        .o_isp6_cis_dvp_h_oe             (o_isp6_cis_dvp_h_oe),
        .o_isp7_cis_dvp_h_oe             (o_isp7_cis_dvp_h_oe),
        .o_isp4_cis_dvp_h_a              (o_isp4_cis_dvp_h_a),
        .o_isp5_cis_dvp_h_a              (o_isp5_cis_dvp_h_a),
        .o_isp6_cis_dvp_h_a              (o_isp6_cis_dvp_h_a),
        .o_isp7_cis_dvp_h_a              (o_isp7_cis_dvp_h_a),
        .o_isp4_cis_dvp_v_oe             (o_isp4_cis_dvp_v_oe),
        .o_isp5_cis_dvp_v_oe             (o_isp5_cis_dvp_v_oe),
        .o_isp6_cis_dvp_v_oe             (o_isp6_cis_dvp_v_oe),
        .o_isp7_cis_dvp_v_oe             (o_isp7_cis_dvp_v_oe),
        .o_isp4_cis_dvp_v_a              (o_isp4_cis_dvp_v_a),
        .o_isp5_cis_dvp_v_a              (o_isp5_cis_dvp_v_a),
        .o_isp6_cis_dvp_v_a              (o_isp6_cis_dvp_v_a),
        .o_isp7_cis_dvp_v_a              (o_isp7_cis_dvp_v_a),
        .MIPI_CLKP_RX4                   (MIPI_CLKP_RX4),
        .MIPI_CLKN_RX4                   (MIPI_CLKN_RX4),
        .MIPI_DP_RX4                     (MIPI_DP_RX4),
        .MIPI_DN_RX4                     (MIPI_DN_RX4),
        .MIPI_CLKP_RX5                   (MIPI_CLKP_RX5),
        .MIPI_CLKN_RX5                   (MIPI_CLKN_RX5),
        .MIPI_DP_RX5                     (MIPI_DP_RX5),
        .MIPI_DN_RX5                     (MIPI_DN_RX5),
        .MIPI_CLKP_RX6                   (MIPI_CLKP_RX6),
        .MIPI_CLKN_RX6                   (MIPI_CLKN_RX6),
        .MIPI_DP_RX6                     (MIPI_DP_RX6),
        .MIPI_DN_RX6                     (MIPI_DN_RX6),
        .MIPI_CLKP_RX7                   (MIPI_CLKP_RX7),
        .MIPI_CLKN_RX7                   (MIPI_CLKN_RX7),
        .MIPI_DP_RX7                     (MIPI_DP_RX7),
        .MIPI_DN_RX7                     (MIPI_DN_RX7),
        .MIPI_CHIP_EN_MR1                (MIPI_CHIP_EN_MR1),
        .MIPI_HS_CKO_RX4                 (MIPI_HS_CKO_RX4),
        .MIPI_HS_DO_RX4                  (MIPI_HS_DO_RX4),
        .MIPI_TEST_VMON_OUT_RX4          (MIPI_TEST_VMON_OUT_RX4),
        .t_aclk                          (t_aclk),
        .t_arstn                         (t_arstn),
        .t_i2cs_scl                      (t_i2cs_scl),
        .t_i_i2cs_sda                    (t_i_i2cs_sda),
        .t_o_i2cs_sda                    (t_o_i2cs_sda),
        .t_isp4_dvp_clk                  (t_isp4_dvp_clk),
        .t_isp4_dvp_v                    (t_isp4_dvp_v),
        .t_isp4_dvp_h                    (t_isp4_dvp_h),
        .t_isp4_dvp_p                    (t_isp4_dvp_p),
        .i_TM_7_MIPI_TEST                (i_TM_7_MIPI_TEST),
        .t_mipi_rx_test_sel              (t_mipi_rx_test_sel),
        .t_clk_isp4                      (t_clk_isp4),
        .t_clk_isp5                      (t_clk_isp5),
        .t_clk_isp6                      (t_clk_isp6),
        .t_clk_isp7                      (t_clk_isp7),
        .t_rstn_isp4                     (t_rstn_isp4),
        .o_fcon_fstart4                  (o_pix4_fstart),
        .o_fcon_fstart5                  (o_pix5_fstart),
        .o_fcon_fstart6                  (o_pix6_fstart),
        .o_fcon_fstart7                  (o_pix7_fstart),
        .i_fcon_mask4                    (i_pix4_mask),
        .i_fcon_mask5                    (i_pix5_mask),
        .i_fcon_mask6                    (i_pix6_mask),
        .i_fcon_mask7                    (i_pix7_mask),
        .o_awuser_isp2main_1             (o_awuser_isp2main_1),
        .o_aruser_isp2main_1             (o_aruser_isp2main_1)
    );

endmodule