//==============================================================================
//
// Project : MVP
//
// Verilog RTL(Behavioral) model
//
// This confidential and proprietary source code may be used only as authorized
// by a licensing agreement from ALPHAHOLDINGS Limited. The entire notice above
// must be reproduced on all authorized copies and copies may only be made to
// the extent permitted by a licensing agreement from ALPHAHOLDINGS Limited.
//
// COPYRIGHT (C) ALPHAHOLDINGS, inc. 2022
//
//==============================================================================
// File name : peri_hpdf
// Version : v1.1
// Description :
// Simulator : NC Verilog
// Created by : bhoh
// Date : 2023-11-15  17:11
//==============================================================================

module peri_hpdf (
    input   [  4:  0]  i_awid_cpu2peri_s0,
    input   [ 31:  0]  i_awaddr_cpu2peri_s0,
    input   [  7:  0]  i_awlen_cpu2peri_s0,
    input   [  2:  0]  i_awsize_cpu2peri_s0,
    input   [  1:  0]  i_awburst_cpu2peri_s0,
    input              i_awlock_cpu2peri_s0,
    input   [  3:  0]  i_awcache_cpu2peri_s0,
    input   [  2:  0]  i_awprot_cpu2peri_s0,
    input              i_awvalid_cpu2peri_s0,
    output             o_awready_cpu2peri_s0,
    input   [ 31:  0]  i_wdata_cpu2peri_s0,
    input   [  3:  0]  i_wstrb_cpu2peri_s0,
    input              i_wlast_cpu2peri_s0,
    input              i_wvalid_cpu2peri_s0,
    output             o_wready_cpu2peri_s0,
    output  [  4:  0]  o_bid_cpu2peri_s0,
    output  [  1:  0]  o_bresp_cpu2peri_s0,
    output             o_bvalid_cpu2peri_s0,
    input              i_bready_cpu2peri_s0,
    input   [  4:  0]  i_arid_cpu2peri_s0,
    input   [ 31:  0]  i_araddr_cpu2peri_s0,
    input   [  7:  0]  i_arlen_cpu2peri_s0,
    input   [  2:  0]  i_arsize_cpu2peri_s0,
    input   [  1:  0]  i_arburst_cpu2peri_s0,
    input              i_arlock_cpu2peri_s0,
    input   [  3:  0]  i_arcache_cpu2peri_s0,
    input   [  2:  0]  i_arprot_cpu2peri_s0,
    input              i_arvalid_cpu2peri_s0,
    output             o_arready_cpu2peri_s0,
    output  [  4:  0]  o_rid_cpu2peri_s0,
    output  [ 31:  0]  o_rdata_cpu2peri_s0,
    output  [  1:  0]  o_rresp_cpu2peri_s0,
    output             o_rlast_cpu2peri_s0,
    output             o_rvalid_cpu2peri_s0,
    input              i_rready_cpu2peri_s0,
    output  [ 31:  0]  o_paddr_peri2ddr_m1,
    output             o_pselx_peri2ddr_m1,
    output             o_penable_peri2ddr_m1,
    output             o_pwrite_peri2ddr_m1,
    input   [ 31:  0]  i_prdata_peri2ddr_m1,
    output  [ 31:  0]  o_pwdata_peri2ddr_m1,
    input              i_pready_peri2ddr_m1,
    input              i_pslverr_peri2ddr_m1,
    output  [ 31:  0]  o_paddr_peri2hsp_m4,
    output             o_pselx_peri2hsp_m4,
    output             o_penable_peri2hsp_m4,
    output             o_pwrite_peri2hsp_m4,
    input   [ 31:  0]  i_prdata_peri2hsp_m4,
    output  [ 31:  0]  o_pwdata_peri2hsp_m4,
    input              i_pready_peri2hsp_m4,
    input              i_pslverr_peri2hsp_m4,
    output  [ 31:  0]  o_paddr_peri2keti_m3,
    output             o_pselx_peri2keti_m3,
    output             o_penable_peri2keti_m3,
    output             o_pwrite_peri2keti_m3,
    input   [ 31:  0]  i_prdata_peri2keti_m3,
    output  [ 31:  0]  o_pwdata_peri2keti_m3,
    input              i_pready_peri2keti_m3,
    input              i_pslverr_peri2keti_m3,
    output  [ 31:  0]  o_haddr_peri2main_m5,
    output  [  2:  0]  o_hburst_peri2main_m5,
    output  [  3:  0]  o_hprot_peri2main_m5,
    output  [  2:  0]  o_hsize_peri2main_m5,
    output  [  1:  0]  o_htrans_peri2main_m5,
    output  [ 31:  0]  o_hwdata_peri2main_m5,
    output             o_hwrite_peri2main_m5,
    input   [ 31:  0]  i_hrdata_peri2main_m5,
    input              i_hresp_peri2main_m5,
    input              i_hready_peri2main_m5,
    output  [ 31:  0]  o_paddr_peri2mna_m2,
    output             o_pselx_peri2mna_m2,
    output             o_penable_peri2mna_m2,
    output             o_pwrite_peri2mna_m2,
    input   [ 31:  0]  i_prdata_peri2mna_m2,
    output  [ 31:  0]  o_pwdata_peri2mna_m2,
    input              i_pready_peri2mna_m2,
    input              i_pslverr_peri2mna_m2,
    input              i_test_bypass,
    input              i_rstn_cpu2peri,
    input              i_clk_cpu2peri,
    input              i_scan_clk,
    input              i_scan_mode,
    input              i_test_rstn,
    output             o_irq_wdt,
    output             o_wdt_nresetout,
    output  [  4:  0]  o_timer0_a,
    output             o_irq_timer0_0,
    output             o_irq_timer0_1,
    output             o_irq_timer0_2,
    output             o_irq_timer0_3,
    output             o_irq_timer0_4,
    output  [  4:  0]  o_timer1_a,
    output             o_irq_timer1_0,
    output             o_irq_timer1_1,
    output             o_irq_timer1_2,
    output             o_irq_timer1_3,
    output             o_irq_timer1_4,
    output             o_irq_uart0,
    input              i_uart0_rxd_y,
    output             o_uart0_txd_a,
    output             o_irq_uart1,
    input              i_uart1_rxd_y,
    output             o_uart1_txd_a,
    input              i_i2c0_scl_y,
    output             o_i2c0_scl_a,
    output             o_i2c0_scl_oe,
    input              i_i2c0_sda_y,
    output             o_i2c0_sda_a,
    output             o_i2c0_sda_oe,
    output             o_irq_i2c0,
    input              i_i2c1_scl_y,
    output             o_i2c1_scl_a,
    output             o_i2c1_scl_oe,
    input              i_i2c1_sda_y,
    output             o_i2c1_sda_a,
    output             o_i2c1_sda_oe,
    output             o_irq_i2c1,
    input              i_i2c2_scl_y,
    output             o_i2c2_scl_a,
    output             o_i2c2_scl_oe,
    input              i_i2c2_sda_y,
    output             o_i2c2_sda_a,
    output             o_i2c2_sda_oe,
    output             o_irq_i2c2,
    input              i_i2c3_scl_y,
    output             o_i2c3_scl_a,
    output             o_i2c3_scl_oe,
    input              i_i2c3_sda_y,
    output             o_i2c3_sda_a,
    output             o_i2c3_sda_oe,
    output             o_irq_i2c3,
    input              i_i2c4_scl_y,
    output             o_i2c4_scl_a,
    output             o_i2c4_scl_oe,
    input              i_i2c4_sda_y,
    output             o_i2c4_sda_a,
    output             o_i2c4_sda_oe,
    output             o_irq_i2c4,
    input              i_i2c5_scl_y,
    output             o_i2c5_scl_a,
    output             o_i2c5_scl_oe,
    input              i_i2c5_sda_y,
    output             o_i2c5_sda_a,
    output             o_i2c5_sda_oe,
    output             o_irq_i2c5,
    input              i_i2c6_scl_y,
    output             o_i2c6_scl_a,
    output             o_i2c6_scl_oe,
    input              i_i2c6_sda_y,
    output             o_i2c6_sda_a,
    output             o_i2c6_sda_oe,
    output             o_irq_i2c6,
    input              i_i2c7_scl_y,
    output             o_i2c7_scl_a,
    output             o_i2c7_scl_oe,
    input              i_i2c7_sda_y,
    output             o_i2c7_sda_a,
    output             o_i2c7_sda_oe,
    output             o_irq_i2c7,
    input              i_i2c8_scl_y,
    output             o_i2c8_scl_a,
    output             o_i2c8_scl_oe,
    input              i_i2c8_sda_y,
    output             o_i2c8_sda_a,
    output             o_i2c8_sda_oe,
    output             o_irq_i2c8,
    input              i_i2c9_scl_y,
    output             o_i2c9_scl_a,
    output             o_i2c9_scl_oe,
    input              i_i2c9_sda_y,
    output             o_i2c9_sda_a,
    output             o_i2c9_sda_oe,
    output             o_irq_i2c9,
    output             o_irq_ssp0,
    output             o_irq_ssp0_txintr,
    output             o_irq_ssp0_rxintr,
    output             o_irq_ssp0_rorintr,
    output             o_irq_ssp0_rtintr,
    input              i_ssp0_clk_y,
    output             o_ssp0_clk_a,
    output             o_ssp0_clk_oe,
    input              i_ssp0_csn_y,
    output             o_ssp0_csn_a,
    output             o_ssp0_csn_oe,
    input              i_ssp0_rx_y,
    output             o_ssp0_tx_a,
    output             o_irq_ssp1,
    output             o_irq_ssp1_txintr,
    output             o_irq_ssp1_rxintr,
    output             o_irq_ssp1_rorintr,
    output             o_irq_ssp1_rtintr,
    input              i_ssp1_clk_y,
    output             o_ssp1_clk_a,
    output             o_ssp1_clk_oe,
    input              i_ssp1_csn_y,
    output             o_ssp1_csn_a,
    output             o_ssp1_csn_oe,
    input              i_ssp1_rx_y,
    output             o_ssp1_tx_a,
    output             o_irq_ssp2,
    output             o_irq_ssp2_txintr,
    output             o_irq_ssp2_rxintr,
    output             o_irq_ssp2_rorintr,
    output             o_irq_ssp2_rtintr,
    input              i_ssp2_clk_y,
    output             o_ssp2_clk_a,
    output             o_ssp2_clk_oe,
    input              i_ssp2_csn_y,
    output             o_ssp2_csn_a,
    output             o_ssp2_csn_oe,
    input              i_ssp2_rx_y,
    output             o_ssp2_tx_a,
    output             o_irq_gpio0,
    input   [  7:  0]  i_gpio0_y,
    output  [  7:  0]  o_gpio0_a,
    output  [  7:  0]  o_gpio0_oe,
    output             o_irq_gpio1,
    input   [  7:  0]  i_gpio1_y,
    output  [  7:  0]  o_gpio1_a,
    output  [  7:  0]  o_gpio1_oe,
    output             o_irq_gpio2,
    input   [  7:  0]  i_gpio2_y,
    output  [  7:  0]  o_gpio2_a,
    output  [  7:  0]  o_gpio2_oe,
    output             o_irq_gpio3,
    input   [  7:  0]  i_gpio3_y,
    output  [  7:  0]  o_gpio3_a,
    output  [  7:  0]  o_gpio3_oe,
    output             o_irq_gpio4,
    input   [  7:  0]  i_gpio4_y,
    output  [  7:  0]  o_gpio4_a,
    output  [  7:  0]  o_gpio4_oe,
    output             o_irq_gpio5,
    input   [  7:  0]  i_gpio5_y,
    output  [  7:  0]  o_gpio5_a,
    output  [  7:  0]  o_gpio5_oe,
    output             o_irq_gpio6,
    input   [  7:  0]  i_gpio6_y,
    output  [  7:  0]  o_gpio6_a,
    output  [  7:  0]  o_gpio6_oe,
    output             o_irq_gpio7,
    input   [  7:  0]  i_gpio7_y,
    output  [  7:  0]  o_gpio7_a,
    output  [  7:  0]  o_gpio7_oe,
    output  [ 19:  0]  o_dmac_breq,
    output  [ 19:  0]  o_dmac_sreq,
    output  [ 19:  0]  o_dmac_lbreq,
    output  [ 19:  0]  o_dmac_lsreq,
    input   [ 19:  0]  i_dmac_clr,
    input   [ 19:  0]  i_dmac_tc,
    input              i_test_mode
);

    wire    [31:0]  peri_bus_paddr_peri_peri0_m0;
    wire            peri_bus_pselx_peri_peri0_m0;
    wire            peri_bus_penable_peri_peri0_m0;
    wire            peri_bus_pwrite_peri_peri0_m0;
    wire    [31:0]  peri_bus_prdata_peri_peri0_m0;
    wire    [31:0]  peri_bus_pwdata_peri_peri0_m0;
    wire            peri_bus_pready_peri_peri0_m0;
    wire            peri_bus_pslverr_peri_peri0_m0;
    wire            peri_crm_o_clk_peri_bus;
    wire            peri_crm_o_rstn_peri_bus;
    wire            peri_crm_o_clk_bus_m0;
    wire            peri_crm_o_rstn_bus_m0;
    wire            peri_crm_o_clk_gpio0;
    wire            peri_crm_o_rstn_gpio0;
    wire            peri_crm_o_clk_gpio1;
    wire            peri_crm_o_rstn_gpio1;
    wire            peri_crm_o_clk_gpio2;
    wire            peri_crm_o_rstn_gpio2;
    wire            peri_crm_o_clk_gpio3;
    wire            peri_crm_o_rstn_gpio3;
    wire            peri_crm_o_clk_gpio4;
    wire            peri_crm_o_rstn_gpio4;
    wire            peri_crm_o_clk_gpio5;
    wire            peri_crm_o_rstn_gpio5;
    wire            peri_crm_o_clk_gpio6;
    wire            peri_crm_o_rstn_gpio6;
    wire            peri_crm_o_clk_gpio7;
    wire            peri_crm_o_rstn_gpio7;
    wire            peri_crm_o_clk_ssp0;
    wire            peri_crm_o_rstn_ssp0;
    wire            peri_crm_o_clk_ssp1;
    wire            peri_crm_o_rstn_ssp1;
    wire            peri_crm_o_clk_ssp2;
    wire            peri_crm_o_rstn_ssp2;
    wire            peri_crm_o_clk_i2c0;
    wire            peri_crm_o_rstn_i2c0;
    wire            peri_crm_o_clk_i2c1;
    wire            peri_crm_o_rstn_i2c1;
    wire            peri_crm_o_clk_i2c2;
    wire            peri_crm_o_rstn_i2c2;
    wire            peri_crm_o_clk_i2c3;
    wire            peri_crm_o_rstn_i2c3;
    wire            peri_crm_o_clk_i2c4;
    wire            peri_crm_o_rstn_i2c4;
    wire            peri_crm_o_clk_i2c5;
    wire            peri_crm_o_rstn_i2c5;
    wire            peri_crm_o_clk_i2c6;
    wire            peri_crm_o_rstn_i2c6;
    wire            peri_crm_o_clk_i2c7;
    wire            peri_crm_o_rstn_i2c7;
    wire            peri_crm_o_clk_i2c8;
    wire            peri_crm_o_rstn_i2c8;
    wire            peri_crm_o_clk_i2c9;
    wire            peri_crm_o_rstn_i2c9;
    wire            peri_crm_o_clk_timer0;
    wire            peri_crm_o_rstn_timer0;
    wire            peri_crm_o_clk_timer1;
    wire            peri_crm_o_rstn_timer1;
    wire            peri_crm_o_clk_uart0;
    wire            peri_crm_o_rstn_uart0;
    wire            peri_crm_o_clk_uart1;
    wire            peri_crm_o_rstn_uart1;
    wire            peri_crm_o_clk_wdt;
    wire            peri_crm_o_rstn_wdt;
    wire            peri_sub_o_crm_apb_psel;
    wire            peri_sub_o_crm_apb_penable;
    wire            peri_sub_o_crm_apb_pwrite;
    wire    [11:0]  peri_sub_o_crm_apb_paddr;
    wire    [31:0]  peri_sub_o_crm_apb_pwdata;
    wire    [31:0]  peri_sub_i_crm_apb_prdata;


    nic400_peri_bus_r0p05 u_peri_bus (
        .awid_cpu2peri_s0        (i_awid_cpu2peri_s0),
        .awaddr_cpu2peri_s0      (i_awaddr_cpu2peri_s0),
        .awlen_cpu2peri_s0       (i_awlen_cpu2peri_s0),
        .awsize_cpu2peri_s0      (i_awsize_cpu2peri_s0),
        .awburst_cpu2peri_s0     (i_awburst_cpu2peri_s0),
        .awlock_cpu2peri_s0      (i_awlock_cpu2peri_s0),
        .awcache_cpu2peri_s0     (i_awcache_cpu2peri_s0),
        .awprot_cpu2peri_s0      (i_awprot_cpu2peri_s0),
        .awvalid_cpu2peri_s0     (i_awvalid_cpu2peri_s0),
        .awready_cpu2peri_s0     (o_awready_cpu2peri_s0),
        .wdata_cpu2peri_s0       (i_wdata_cpu2peri_s0),
        .wstrb_cpu2peri_s0       (i_wstrb_cpu2peri_s0),
        .wlast_cpu2peri_s0       (i_wlast_cpu2peri_s0),
        .wvalid_cpu2peri_s0      (i_wvalid_cpu2peri_s0),
        .wready_cpu2peri_s0      (o_wready_cpu2peri_s0),
        .bid_cpu2peri_s0         (o_bid_cpu2peri_s0),
        .bresp_cpu2peri_s0       (o_bresp_cpu2peri_s0),
        .bvalid_cpu2peri_s0      (o_bvalid_cpu2peri_s0),
        .bready_cpu2peri_s0      (i_bready_cpu2peri_s0),
        .arid_cpu2peri_s0        (i_arid_cpu2peri_s0),
        .araddr_cpu2peri_s0      (i_araddr_cpu2peri_s0),
        .arlen_cpu2peri_s0       (i_arlen_cpu2peri_s0),
        .arsize_cpu2peri_s0      (i_arsize_cpu2peri_s0),
        .arburst_cpu2peri_s0     (i_arburst_cpu2peri_s0),
        .arlock_cpu2peri_s0      (i_arlock_cpu2peri_s0),
        .arcache_cpu2peri_s0     (i_arcache_cpu2peri_s0),
        .arprot_cpu2peri_s0      (i_arprot_cpu2peri_s0),
        .arvalid_cpu2peri_s0     (i_arvalid_cpu2peri_s0),
        .arready_cpu2peri_s0     (o_arready_cpu2peri_s0),
        .rid_cpu2peri_s0         (o_rid_cpu2peri_s0),
        .rdata_cpu2peri_s0       (o_rdata_cpu2peri_s0),
        .rresp_cpu2peri_s0       (o_rresp_cpu2peri_s0),
        .rlast_cpu2peri_s0       (o_rlast_cpu2peri_s0),
        .rvalid_cpu2peri_s0      (o_rvalid_cpu2peri_s0),
        .rready_cpu2peri_s0      (i_rready_cpu2peri_s0),
        .paddr_peri2ddr_m1       (o_paddr_peri2ddr_m1),
        .pselx_peri2ddr_m1       (o_pselx_peri2ddr_m1),
        .penable_peri2ddr_m1     (o_penable_peri2ddr_m1),
        .pwrite_peri2ddr_m1      (o_pwrite_peri2ddr_m1),
        .prdata_peri2ddr_m1      (i_prdata_peri2ddr_m1),
        .pwdata_peri2ddr_m1      (o_pwdata_peri2ddr_m1),
        .pready_peri2ddr_m1      (i_pready_peri2ddr_m1),
        .pslverr_peri2ddr_m1     (i_pslverr_peri2ddr_m1),
        .paddr_peri2hsp_m4       (o_paddr_peri2hsp_m4),
        .pselx_peri2hsp_m4       (o_pselx_peri2hsp_m4),
        .penable_peri2hsp_m4     (o_penable_peri2hsp_m4),
        .pwrite_peri2hsp_m4      (o_pwrite_peri2hsp_m4),
        .prdata_peri2hsp_m4      (i_prdata_peri2hsp_m4),
        .pwdata_peri2hsp_m4      (o_pwdata_peri2hsp_m4),
        .pready_peri2hsp_m4      (i_pready_peri2hsp_m4),
        .pslverr_peri2hsp_m4     (i_pslverr_peri2hsp_m4),
        .paddr_peri2keti_m3      (o_paddr_peri2keti_m3),
        .pselx_peri2keti_m3      (o_pselx_peri2keti_m3),
        .penable_peri2keti_m3    (o_penable_peri2keti_m3),
        .pwrite_peri2keti_m3     (o_pwrite_peri2keti_m3),
        .prdata_peri2keti_m3     (i_prdata_peri2keti_m3),
        .pwdata_peri2keti_m3     (o_pwdata_peri2keti_m3),
        .pready_peri2keti_m3     (i_pready_peri2keti_m3),
        .pslverr_peri2keti_m3    (i_pslverr_peri2keti_m3),
        .haddr_peri2main_m5      (o_haddr_peri2main_m5),
        .hburst_peri2main_m5     (o_hburst_peri2main_m5),
        .hprot_peri2main_m5      (o_hprot_peri2main_m5),
        .hsize_peri2main_m5      (o_hsize_peri2main_m5),
        .htrans_peri2main_m5     (o_htrans_peri2main_m5),
        .hwdata_peri2main_m5     (o_hwdata_peri2main_m5),
        .hwrite_peri2main_m5     (o_hwrite_peri2main_m5),
        .hrdata_peri2main_m5     (i_hrdata_peri2main_m5),
        .hresp_peri2main_m5      (i_hresp_peri2main_m5),
        .hready_peri2main_m5     (i_hready_peri2main_m5),
        .paddr_peri2mna_m2       (o_paddr_peri2mna_m2),
        .pselx_peri2mna_m2       (o_pselx_peri2mna_m2),
        .penable_peri2mna_m2     (o_penable_peri2mna_m2),
        .pwrite_peri2mna_m2      (o_pwrite_peri2mna_m2),
        .prdata_peri2mna_m2      (i_prdata_peri2mna_m2),
        .pwdata_peri2mna_m2      (o_pwdata_peri2mna_m2),
        .pready_peri2mna_m2      (i_pready_peri2mna_m2),
        .pslverr_peri2mna_m2     (i_pslverr_peri2mna_m2),
        .paddr_peri_peri0_m0     (peri_bus_paddr_peri_peri0_m0),
        .pselx_peri_peri0_m0     (peri_bus_pselx_peri_peri0_m0),
        .penable_peri_peri0_m0   (peri_bus_penable_peri_peri0_m0),
        .pwrite_peri_peri0_m0    (peri_bus_pwrite_peri_peri0_m0),
        .prdata_peri_peri0_m0    (peri_bus_prdata_peri_peri0_m0),
        .pwdata_peri_peri0_m0    (peri_bus_pwdata_peri_peri0_m0),
        .pready_peri_peri0_m0    (peri_bus_pready_peri_peri0_m0),
        .pslverr_peri_peri0_m0   (peri_bus_pslverr_peri_peri0_m0),
        .mainclk                 (peri_crm_o_clk_peri_bus),
        .mainclk_r               (peri_crm_o_clk_peri_bus),
        .mainclken               (1'h1),
        .mainresetn              (peri_crm_o_rstn_peri_bus),
        .mainresetn_r            (peri_crm_o_rstn_peri_bus)
    );

    mvp_crm_peri u_peri_crm (
        .i_test_bypass           (i_test_bypass),
        .i_rstn_peri             (i_rstn_cpu2peri),
        .i_apb_pclk              (i_clk_cpu2peri),
        .i_apb_prstn             (i_rstn_cpu2peri),
        .i_apb_psel              (peri_sub_o_crm_apb_psel),
        .i_apb_penable           (peri_sub_o_crm_apb_penable),
        .i_apb_pwrite            (peri_sub_o_crm_apb_pwrite),
        .i_apb_paddr             (peri_sub_o_crm_apb_paddr),
        .i_apb_pwdata            (peri_sub_o_crm_apb_pwdata),
        .o_apb_prdata            (peri_sub_i_crm_apb_prdata),
        .i_clk_cpu2peri          (i_clk_cpu2peri),
        .o_clk_peri_bus          (peri_crm_o_clk_peri_bus),
        .o_rstn_peri_bus         (peri_crm_o_rstn_peri_bus),
        .o_clk_bus_m0            (peri_crm_o_clk_bus_m0),
        .o_rstn_bus_m0           (peri_crm_o_rstn_bus_m0),
        .o_clk_gpio0             (peri_crm_o_clk_gpio0),
        .o_rstn_gpio0            (peri_crm_o_rstn_gpio0),
        .o_clk_gpio1             (peri_crm_o_clk_gpio1),
        .o_rstn_gpio1            (peri_crm_o_rstn_gpio1),
        .o_clk_gpio2             (peri_crm_o_clk_gpio2),
        .o_rstn_gpio2            (peri_crm_o_rstn_gpio2),
        .o_clk_gpio3             (peri_crm_o_clk_gpio3),
        .o_rstn_gpio3            (peri_crm_o_rstn_gpio3),
        .o_clk_gpio4             (peri_crm_o_clk_gpio4),
        .o_rstn_gpio4            (peri_crm_o_rstn_gpio4),
        .o_clk_gpio5             (peri_crm_o_clk_gpio5),
        .o_rstn_gpio5            (peri_crm_o_rstn_gpio5),
        .o_clk_gpio6             (peri_crm_o_clk_gpio6),
        .o_rstn_gpio6            (peri_crm_o_rstn_gpio6),
        .o_clk_gpio7             (peri_crm_o_clk_gpio7),
        .o_rstn_gpio7            (peri_crm_o_rstn_gpio7),
        .o_clk_ssp0              (peri_crm_o_clk_ssp0),
        .o_rstn_ssp0             (peri_crm_o_rstn_ssp0),
        .o_clk_ssp1              (peri_crm_o_clk_ssp1),
        .o_rstn_ssp1             (peri_crm_o_rstn_ssp1),
        .o_clk_ssp2              (peri_crm_o_clk_ssp2),
        .o_rstn_ssp2             (peri_crm_o_rstn_ssp2),
        .o_clk_i2c0              (peri_crm_o_clk_i2c0),
        .o_rstn_i2c0             (peri_crm_o_rstn_i2c0),
        .o_clk_i2c1              (peri_crm_o_clk_i2c1),
        .o_rstn_i2c1             (peri_crm_o_rstn_i2c1),
        .o_clk_i2c2              (peri_crm_o_clk_i2c2),
        .o_rstn_i2c2             (peri_crm_o_rstn_i2c2),
        .o_clk_i2c3              (peri_crm_o_clk_i2c3),
        .o_rstn_i2c3             (peri_crm_o_rstn_i2c3),
        .o_clk_i2c4              (peri_crm_o_clk_i2c4),
        .o_rstn_i2c4             (peri_crm_o_rstn_i2c4),
        .o_clk_i2c5              (peri_crm_o_clk_i2c5),
        .o_rstn_i2c5             (peri_crm_o_rstn_i2c5),
        .o_clk_i2c6              (peri_crm_o_clk_i2c6),
        .o_rstn_i2c6             (peri_crm_o_rstn_i2c6),
        .o_clk_i2c7              (peri_crm_o_clk_i2c7),
        .o_rstn_i2c7             (peri_crm_o_rstn_i2c7),
        .o_clk_i2c8              (peri_crm_o_clk_i2c8),
        .o_rstn_i2c8             (peri_crm_o_rstn_i2c8),
        .o_clk_i2c9              (peri_crm_o_clk_i2c9),
        .o_rstn_i2c9             (peri_crm_o_rstn_i2c9),
        .o_clk_timer0            (peri_crm_o_clk_timer0),
        .o_rstn_timer0           (peri_crm_o_rstn_timer0),
        .o_clk_timer1            (peri_crm_o_clk_timer1),
        .o_rstn_timer1           (peri_crm_o_rstn_timer1),
        .o_clk_uart0             (peri_crm_o_clk_uart0),
        .o_rstn_uart0            (peri_crm_o_rstn_uart0),
        .o_clk_uart1             (peri_crm_o_clk_uart1),
        .o_rstn_uart1            (peri_crm_o_rstn_uart1),
        .o_clk_wdt               (peri_crm_o_clk_wdt),
        .o_rstn_wdt              (peri_crm_o_rstn_wdt),
        .i_scan_clk              (i_scan_clk),
        .i_scan_mode             (i_scan_mode),
        .i_scan_rstn             (i_test_rstn)
    );

    peri_sub u_peri_sub (
        .i_clk_bus_m0            (peri_crm_o_clk_bus_m0),
        .i_rstn_bus_m0           (peri_crm_o_rstn_bus_m0),
        .i_clk_gpio0             (peri_crm_o_clk_gpio0),
        .i_rstn_gpio0            (peri_crm_o_rstn_gpio0),
        .i_clk_gpio1             (peri_crm_o_clk_gpio1),
        .i_rstn_gpio1            (peri_crm_o_rstn_gpio1),
        .i_clk_gpio2             (peri_crm_o_clk_gpio2),
        .i_rstn_gpio2            (peri_crm_o_rstn_gpio2),
        .i_clk_gpio3             (peri_crm_o_clk_gpio3),
        .i_rstn_gpio3            (peri_crm_o_rstn_gpio3),
        .i_clk_gpio4             (peri_crm_o_clk_gpio4),
        .i_rstn_gpio4            (peri_crm_o_rstn_gpio4),
        .i_clk_gpio5             (peri_crm_o_clk_gpio5),
        .i_rstn_gpio5            (peri_crm_o_rstn_gpio5),
        .i_clk_gpio6             (peri_crm_o_clk_gpio6),
        .i_rstn_gpio6            (peri_crm_o_rstn_gpio6),
        .i_clk_gpio7             (peri_crm_o_clk_gpio7),
        .i_rstn_gpio7            (peri_crm_o_rstn_gpio7),
        .i_clk_ssp0              (peri_crm_o_clk_ssp0),
        .i_rstn_ssp0             (peri_crm_o_rstn_ssp0),
        .i_clk_ssp1              (peri_crm_o_clk_ssp1),
        .i_rstn_ssp1             (peri_crm_o_rstn_ssp1),
        .i_clk_ssp2              (peri_crm_o_clk_ssp2),
        .i_rstn_ssp2             (peri_crm_o_rstn_ssp2),
        .i_clk_i2c0              (peri_crm_o_clk_i2c0),
        .i_rstn_i2c0             (peri_crm_o_rstn_i2c0),
        .i_clk_i2c1              (peri_crm_o_clk_i2c1),
        .i_rstn_i2c1             (peri_crm_o_rstn_i2c1),
        .i_clk_i2c2              (peri_crm_o_clk_i2c2),
        .i_rstn_i2c2             (peri_crm_o_rstn_i2c2),
        .i_clk_i2c3              (peri_crm_o_clk_i2c3),
        .i_rstn_i2c3             (peri_crm_o_rstn_i2c3),
        .i_clk_i2c4              (peri_crm_o_clk_i2c4),
        .i_rstn_i2c4             (peri_crm_o_rstn_i2c4),
        .i_clk_i2c5              (peri_crm_o_clk_i2c5),
        .i_rstn_i2c5             (peri_crm_o_rstn_i2c5),
        .i_clk_i2c6              (peri_crm_o_clk_i2c6),
        .i_rstn_i2c6             (peri_crm_o_rstn_i2c6),
        .i_clk_i2c7              (peri_crm_o_clk_i2c7),
        .i_rstn_i2c7             (peri_crm_o_rstn_i2c7),
        .i_clk_i2c8              (peri_crm_o_clk_i2c8),
        .i_rstn_i2c8             (peri_crm_o_rstn_i2c8),
        .i_clk_i2c9              (peri_crm_o_clk_i2c9),
        .i_rstn_i2c9             (peri_crm_o_rstn_i2c9),
        .i_clk_pwm0              (peri_crm_o_clk_timer0),
        .i_rstn_pwm0             (peri_crm_o_rstn_timer0),
        .i_clk_pwm1              (peri_crm_o_clk_timer1),
        .i_rstn_pwm1             (peri_crm_o_rstn_timer1),
        .i_clk_uart0             (peri_crm_o_clk_uart0),
        .i_rstn_uart0            (peri_crm_o_rstn_uart0),
        .i_clk_uart1             (peri_crm_o_clk_uart1),
        .i_rstn_uart1            (peri_crm_o_rstn_uart1),
        .i_clk_wdt0              (peri_crm_o_clk_wdt),
        .i_rstn_wdt0             (peri_crm_o_rstn_wdt),
        .o_crm_apb_psel          (peri_sub_o_crm_apb_psel),
        .o_crm_apb_penable       (peri_sub_o_crm_apb_penable),
        .o_crm_apb_pwrite        (peri_sub_o_crm_apb_pwrite),
        .o_crm_apb_paddr         (peri_sub_o_crm_apb_paddr),
        .o_crm_apb_pwdata        (peri_sub_o_crm_apb_pwdata),
        .i_crm_apb_prdata        (peri_sub_i_crm_apb_prdata),
        .i_paddr_peri0_m0        (peri_bus_paddr_peri_peri0_m0),
        .i_pselx_peri0_m0        (peri_bus_pselx_peri_peri0_m0),
        .i_penable_peri0_m0      (peri_bus_penable_peri_peri0_m0),
        .i_pwrite_peri0_m0       (peri_bus_pwrite_peri_peri0_m0),
        .o_prdata_peri0_m0       (peri_bus_prdata_peri_peri0_m0),
        .i_pwdata_peri0_m0       (peri_bus_pwdata_peri_peri0_m0),
        .o_pready_peri0_m0       (peri_bus_pready_peri_peri0_m0),
        .o_pslverr_peri0_m0      (peri_bus_pslverr_peri_peri0_m0),
        .o_irq_wdt               (o_irq_wdt),
        .o_wdt_nresetout         (o_wdt_nresetout),
        .o_timer0_a              (o_timer0_a),
        .o_irq_timer0_0          (o_irq_timer0_0),
        .o_irq_timer0_1          (o_irq_timer0_1),
        .o_irq_timer0_2          (o_irq_timer0_2),
        .o_irq_timer0_3          (o_irq_timer0_3),
        .o_irq_timer0_4          (o_irq_timer0_4),
        .o_timer1_a              (o_timer1_a),
        .o_irq_timer1_0          (o_irq_timer1_0),
        .o_irq_timer1_1          (o_irq_timer1_1),
        .o_irq_timer1_2          (o_irq_timer1_2),
        .o_irq_timer1_3          (o_irq_timer1_3),
        .o_irq_timer1_4          (o_irq_timer1_4),
        .o_irq_uart0             (o_irq_uart0),
        .i_uart0_rxd_y           (i_uart0_rxd_y),
        .o_uart0_txd_a           (o_uart0_txd_a),
        .o_irq_uart1             (o_irq_uart1),
        .i_uart1_rxd_y           (i_uart1_rxd_y),
        .o_uart1_txd_a           (o_uart1_txd_a),
        .i_i2c0_scl_y            (i_i2c0_scl_y),
        .o_i2c0_scl_a            (o_i2c0_scl_a),
        .o_i2c0_scl_oe           (o_i2c0_scl_oe),
        .i_i2c0_sda_y            (i_i2c0_sda_y),
        .o_i2c0_sda_a            (o_i2c0_sda_a),
        .o_i2c0_sda_oe           (o_i2c0_sda_oe),
        .o_irq_i2c0              (o_irq_i2c0),
        .i_i2c1_scl_y            (i_i2c1_scl_y),
        .o_i2c1_scl_a            (o_i2c1_scl_a),
        .o_i2c1_scl_oe           (o_i2c1_scl_oe),
        .i_i2c1_sda_y            (i_i2c1_sda_y),
        .o_i2c1_sda_a            (o_i2c1_sda_a),
        .o_i2c1_sda_oe           (o_i2c1_sda_oe),
        .o_irq_i2c1              (o_irq_i2c1),
        .i_i2c2_scl_y            (i_i2c2_scl_y),
        .o_i2c2_scl_a            (o_i2c2_scl_a),
        .o_i2c2_scl_oe           (o_i2c2_scl_oe),
        .i_i2c2_sda_y            (i_i2c2_sda_y),
        .o_i2c2_sda_a            (o_i2c2_sda_a),
        .o_i2c2_sda_oe           (o_i2c2_sda_oe),
        .o_irq_i2c2              (o_irq_i2c2),
        .i_i2c3_scl_y            (i_i2c3_scl_y),
        .o_i2c3_scl_a            (o_i2c3_scl_a),
        .o_i2c3_scl_oe           (o_i2c3_scl_oe),
        .i_i2c3_sda_y            (i_i2c3_sda_y),
        .o_i2c3_sda_a            (o_i2c3_sda_a),
        .o_i2c3_sda_oe           (o_i2c3_sda_oe),
        .o_irq_i2c3              (o_irq_i2c3),
        .i_i2c4_scl_y            (i_i2c4_scl_y),
        .o_i2c4_scl_a            (o_i2c4_scl_a),
        .o_i2c4_scl_oe           (o_i2c4_scl_oe),
        .i_i2c4_sda_y            (i_i2c4_sda_y),
        .o_i2c4_sda_a            (o_i2c4_sda_a),
        .o_i2c4_sda_oe           (o_i2c4_sda_oe),
        .o_irq_i2c4              (o_irq_i2c4),
        .i_i2c5_scl_y            (i_i2c5_scl_y),
        .o_i2c5_scl_a            (o_i2c5_scl_a),
        .o_i2c5_scl_oe           (o_i2c5_scl_oe),
        .i_i2c5_sda_y            (i_i2c5_sda_y),
        .o_i2c5_sda_a            (o_i2c5_sda_a),
        .o_i2c5_sda_oe           (o_i2c5_sda_oe),
        .o_irq_i2c5              (o_irq_i2c5),
        .i_i2c6_scl_y            (i_i2c6_scl_y),
        .o_i2c6_scl_a            (o_i2c6_scl_a),
        .o_i2c6_scl_oe           (o_i2c6_scl_oe),
        .i_i2c6_sda_y            (i_i2c6_sda_y),
        .o_i2c6_sda_a            (o_i2c6_sda_a),
        .o_i2c6_sda_oe           (o_i2c6_sda_oe),
        .o_irq_i2c6              (o_irq_i2c6),
        .i_i2c7_scl_y            (i_i2c7_scl_y),
        .o_i2c7_scl_a            (o_i2c7_scl_a),
        .o_i2c7_scl_oe           (o_i2c7_scl_oe),
        .i_i2c7_sda_y            (i_i2c7_sda_y),
        .o_i2c7_sda_a            (o_i2c7_sda_a),
        .o_i2c7_sda_oe           (o_i2c7_sda_oe),
        .o_irq_i2c7              (o_irq_i2c7),
        .i_i2c8_scl_y            (i_i2c8_scl_y),
        .o_i2c8_scl_a            (o_i2c8_scl_a),
        .o_i2c8_scl_oe           (o_i2c8_scl_oe),
        .i_i2c8_sda_y            (i_i2c8_sda_y),
        .o_i2c8_sda_a            (o_i2c8_sda_a),
        .o_i2c8_sda_oe           (o_i2c8_sda_oe),
        .o_irq_i2c8              (o_irq_i2c8),
        .i_i2c9_scl_y            (i_i2c9_scl_y),
        .o_i2c9_scl_a            (o_i2c9_scl_a),
        .o_i2c9_scl_oe           (o_i2c9_scl_oe),
        .i_i2c9_sda_y            (i_i2c9_sda_y),
        .o_i2c9_sda_a            (o_i2c9_sda_a),
        .o_i2c9_sda_oe           (o_i2c9_sda_oe),
        .o_irq_i2c9              (o_irq_i2c9),
        .o_irq_ssp0              (o_irq_ssp0),
        .o_irq_ssp0_txintr       (o_irq_ssp0_txintr),
        .o_irq_ssp0_rxintr       (o_irq_ssp0_rxintr),
        .o_irq_ssp0_rorintr      (o_irq_ssp0_rorintr),
        .o_irq_ssp0_rtintr       (o_irq_ssp0_rtintr),
        .i_ssp0_clk_y            (i_ssp0_clk_y),
        .o_ssp0_clk_a            (o_ssp0_clk_a),
        .o_ssp0_clk_oe           (o_ssp0_clk_oe),
        .i_ssp0_csn_y            (i_ssp0_csn_y),
        .o_ssp0_csn_a            (o_ssp0_csn_a),
        .o_ssp0_csn_oe           (o_ssp0_csn_oe),
        .i_ssp0_rx_y             (i_ssp0_rx_y),
        .o_ssp0_tx_a             (o_ssp0_tx_a),
        .o_irq_ssp1              (o_irq_ssp1),
        .o_irq_ssp1_txintr       (o_irq_ssp1_txintr),
        .o_irq_ssp1_rxintr       (o_irq_ssp1_rxintr),
        .o_irq_ssp1_rorintr      (o_irq_ssp1_rorintr),
        .o_irq_ssp1_rtintr       (o_irq_ssp1_rtintr),
        .i_ssp1_clk_y            (i_ssp1_clk_y),
        .o_ssp1_clk_a            (o_ssp1_clk_a),
        .o_ssp1_clk_oe           (o_ssp1_clk_oe),
        .i_ssp1_csn_y            (i_ssp1_csn_y),
        .o_ssp1_csn_a            (o_ssp1_csn_a),
        .o_ssp1_csn_oe           (o_ssp1_csn_oe),
        .i_ssp1_rx_y             (i_ssp1_rx_y),
        .o_ssp1_tx_a             (o_ssp1_tx_a),
        .o_irq_ssp2              (o_irq_ssp2),
        .o_irq_ssp2_txintr       (o_irq_ssp2_txintr),
        .o_irq_ssp2_rxintr       (o_irq_ssp2_rxintr),
        .o_irq_ssp2_rorintr      (o_irq_ssp2_rorintr),
        .o_irq_ssp2_rtintr       (o_irq_ssp2_rtintr),
        .i_ssp2_clk_y            (i_ssp2_clk_y),
        .o_ssp2_clk_a            (o_ssp2_clk_a),
        .o_ssp2_clk_oe           (o_ssp2_clk_oe),
        .i_ssp2_csn_y            (i_ssp2_csn_y),
        .o_ssp2_csn_a            (o_ssp2_csn_a),
        .o_ssp2_csn_oe           (o_ssp2_csn_oe),
        .i_ssp2_rx_y             (i_ssp2_rx_y),
        .o_ssp2_tx_a             (o_ssp2_tx_a),
        .o_irq_gpio0             (o_irq_gpio0),
        .i_gpio0_y               (i_gpio0_y),
        .o_gpio0_a               (o_gpio0_a),
        .o_gpio0_oe              (o_gpio0_oe),
        .o_irq_gpio1             (o_irq_gpio1),
        .i_gpio1_y               (i_gpio1_y),
        .o_gpio1_a               (o_gpio1_a),
        .o_gpio1_oe              (o_gpio1_oe),
        .o_irq_gpio2             (o_irq_gpio2),
        .i_gpio2_y               (i_gpio2_y),
        .o_gpio2_a               (o_gpio2_a),
        .o_gpio2_oe              (o_gpio2_oe),
        .o_irq_gpio3             (o_irq_gpio3),
        .i_gpio3_y               (i_gpio3_y),
        .o_gpio3_a               (o_gpio3_a),
        .o_gpio3_oe              (o_gpio3_oe),
        .o_irq_gpio4             (o_irq_gpio4),
        .i_gpio4_y               (i_gpio4_y),
        .o_gpio4_a               (o_gpio4_a),
        .o_gpio4_oe              (o_gpio4_oe),
        .o_irq_gpio5             (o_irq_gpio5),
        .i_gpio5_y               (i_gpio5_y),
        .o_gpio5_a               (o_gpio5_a),
        .o_gpio5_oe              (o_gpio5_oe),
        .o_irq_gpio6             (o_irq_gpio6),
        .i_gpio6_y               (i_gpio6_y),
        .o_gpio6_a               (o_gpio6_a),
        .o_gpio6_oe              (o_gpio6_oe),
        .o_irq_gpio7             (o_irq_gpio7),
        .i_gpio7_y               (i_gpio7_y),
        .o_gpio7_a               (o_gpio7_a),
        .o_gpio7_oe              (o_gpio7_oe),
        .o_dmac_breq             (o_dmac_breq),
        .o_dmac_sreq             (o_dmac_sreq),
        .o_dmac_lbreq            (o_dmac_lbreq),
        .o_dmac_lsreq            (o_dmac_lsreq),
        .i_dmac_clr              (i_dmac_clr),
        .i_dmac_tc               (i_dmac_tc),
        .i_test_mode             (i_test_mode)
    );

endmodule