

module analog_top (
    input   [  1:  0]   i_pll2551_mode,
    input   [  5:  0]   i_norm_p,
    input   [  9:  0]   i_norm_m,
    input   [  2:  0]   i_norm_s,
    input   [  1:  0]   i_norm_lock_con_in,
    input   [  1:  0]   i_norm_lock_con_out,
    input   [  1:  0]   i_norm_lock_con_dly,
    input   [  1:  0]   i_norm_lock_con_rev,
    input   [  4:  0]   i_norm_tst_afc,
    input   [  1:  0]   i_norm_icp,
    input               i_norm_fin,
    input               i_norm_resetb,
    input               i_norm_bypass,
    input               i_norm_tst_en,
    input               i_norm_fsel,
    input               i_norm_feed_en,
    input               i_norm_lock_en,
    input               i_norm_afcini_sel,
    input               i_norm_vcoini_en,
    input               i_norm_fout_mask,
    input               i_norm_pbias_ctrl,
    input               i_norm_pbias_ctrl_en,
    input   [  5:  0]   t_main_pll_p,
    input   [  9:  0]   t_main_pll_m,
    input   [  2:  0]   t_main_pll_s,
    input   [  1:  0]   t_main_pll_lock_con_in,
    input   [  1:  0]   t_main_pll_lock_con_out,
    input   [  1:  0]   t_main_pll_lock_con_dly,
    input   [  1:  0]   t_main_pll_lock_con_rev,
    input   [  4:  0]   t_main_pll_tst_afc,
    input   [  1:  0]   t_main_pll_icp,
    input               t_main_pll_resetb,
    input               t_main_pll_bypass,
    input               t_main_pll_tst_en,
    input               t_main_pll_fsel,
    input               t_main_pll_feed_en,
    input               t_main_pll_lock_en,
    input               t_main_pll_afcini_sel,
    input               t_main_pll_vcoini_en,
    input               t_main_pll_fout_mask,
    input               t_main_pll_pbias_ctrl,
    input               t_main_pll_pbias_ctrl_en,
    output              o_feed_out,
    output              o_lock,
    output              o_fout,
    output              o_sync_m_clk_out,
    output  [  4:  0]   o_afc_code,
    output              t_main_pll_feed_out,
    output              t_main_pll_lock,
    output              t_main_pll_fout,
    output              t_main_pll_sync_m_clk_out,
    output  [  4:  0]   t_main_pll_afc_code,
    input   [  5:  0]   sr_main_pll_p,
    input   [  9:  0]   sr_main_pll_m,
    input   [  2:  0]   sr_main_pll_s,
    output              o_por_sys
); 

    tmux_sf_pll2551x_ln28lpp_5000 u_tmux_sf_pll2551x(
        .i_tmode		        (i_pll2551_mode	        ),
        .i_norm_p		        (i_norm_p		        ),
        .i_norm_m		        (i_norm_m		        ),
        .i_norm_s		        (i_norm_s		        ),
        .i_norm_lock_con_in		(i_norm_lock_con_in	    ),
        .i_norm_lock_con_out    (i_norm_lock_con_out    ),
        .i_norm_lock_con_dly    (i_norm_lock_con_dly    ),
        .i_norm_lock_con_rev    (i_norm_lock_con_rev    ),
        .i_norm_tst_afc		    (i_norm_tst_afc		    ),
        .i_norm_icp		        (i_norm_icp		        ),
        .i_norm_fin		        (i_norm_fin		        ),
        .i_norm_resetb		    (i_norm_resetb		    ),
        .i_norm_bypass		    (i_norm_bypass		    ),
        .i_norm_tst_en		    (i_norm_tst_en		    ),
        .i_norm_fsel		    (i_norm_fsel		    ),
        .i_norm_feed_en		    (i_norm_feed_en		    ),
        .i_norm_lock_en		    (i_norm_lock_en		    ),
        .i_norm_afcini_sel		(i_norm_afcini_sel	    ),
        .i_norm_vcoini_en		(i_norm_vcoini_en	    ),
        .i_norm_fout_mask		(i_norm_fout_mask	    ),
        .i_norm_pbias_ctrl		(i_norm_pbias_ctrl	    ),
        .i_norm_pbias_ctrl_en	(i_norm_pbias_ctrl_en   ),
        .i_test0_p		        (t_main_pll_p               ),
        .i_test0_m		        (t_main_pll_m               ),
        .i_test0_s		        (t_main_pll_s               ),
        .i_test0_lock_con_in	(t_main_pll_lock_con_in     ),
        .i_test0_lock_con_out	(t_main_pll_lock_con_out    ),
        .i_test0_lock_con_dly	(t_main_pll_lock_con_dly    ),
        .i_test0_lock_con_rev	(t_main_pll_lock_con_rev    ),
        .i_test0_tst_afc		(t_main_pll_tst_afc         ),
        .i_test0_icp		    (t_main_pll_icp             ),
        .i_test0_fin		    (i_norm_fin                 ),
        .i_test0_resetb		    (t_main_pll_resetb          ),
        .i_test0_bypass		    (t_main_pll_bypass          ),
        .i_test0_tst_en		    (t_main_pll_tst_en          ),
        .i_test0_fsel		    (t_main_pll_fsel            ),
        .i_test0_feed_en		(t_main_pll_feed_en         ),
        .i_test0_lock_en		(t_main_pll_lock_en         ),
        .i_test0_afcini_sel		(t_main_pll_afcini_sel      ),
        .i_test0_vcoini_en		(t_main_pll_vcoini_en       ),
        .i_test0_fout_mask		(t_main_pll_fout_mask       ),
        .i_test0_pbias_ctrl		(t_main_pll_pbias_ctrl      ),
        .i_test0_pbias_ctrl_en	(t_main_pll_pbias_ctrl_en   ),
        .i_test1_p		        (sr_main_pll_p              ),
        .i_test1_m		        (sr_main_pll_m              ),
        .i_test1_s		        (sr_main_pll_s              ),
        .i_test1_lock_con_in	(2'h3                       ),
        .i_test1_lock_con_out	(2'h3                       ),
        .i_test1_lock_con_dly	(2'h3                       ),
        .i_test1_lock_con_rev	(2'h0                       ),
        .i_test1_tst_afc		(5'h0                       ),
        .i_test1_icp		    (2'h0                       ),
        .i_test1_fin		    (i_norm_fin                 ),
        .i_test1_resetb		    (t_main_pll_resetb          ),
        .i_test1_bypass		    (1'h0                       ),
        .i_test1_tst_en		    (1'h0                       ),
        .i_test1_fsel		    (1'h0                       ),
        .i_test1_feed_en		(1'h0                       ),
        .i_test1_lock_en		(1'h1                       ),
        .i_test1_afcini_sel		(1'h0                       ),
        .i_test1_vcoini_en		(1'h1                       ),
        .i_test1_fout_mask		(1'h0                       ),
        .i_test1_pbias_ctrl		(1'h0                       ),
        .i_test1_pbias_ctrl_en	(1'h0                       ),
        .o_feed_out		        (o_feed_out		            ),
        .o_lock		            (o_lock		                ),
        .o_fout		            (o_fout		                ),
        .o_sync_m_clk_out		(o_sync_m_clk_out		    ),
        .o_afc_code             (o_afc_code                 )
    );

    assign t_main_pll_feed_out		    = o_feed_out;		
    assign t_main_pll_lock		        = o_lock;		
    assign t_main_pll_fout		        = o_fout;		
    assign t_main_pll_sync_m_clk_out    = o_sync_m_clk_out;			
    assign t_main_pll_afc_code		    = o_afc_code;		



    sf_por2803xa_ln28lpp    u_sf_por2803xa_ln28lpp ( 
        .SYS    ( o_por_sys    ) // System Power on Reset for internal
    );

endmodule 
