module slave_axi_128 (
    input           i_aclk    ,
    input           i_aresetn ,
    input  [3:0]    i_awid    ,
    input  [31:0]   i_awaddr  ,
    input  [3:0]    i_awlen   ,
    input  [2:0]    i_awsize  ,
    input  [1:0]    i_awburst ,
    input  [1:0]    i_awlock  ,
    input  [3:0]    i_awcache ,
    input  [2:0]    i_awprot  ,
    input           i_awvalid ,
    output          o_awready ,
    input  [3:0]    i_wid     ,
    input  [127:0]  i_wdata   ,
    input  [15:0]   i_wstrb   ,
    input           i_wlast   ,
    input           i_wvalid  ,
    output          o_wready  ,
    output [3:0]    o_bid     ,
    output [1:0]    o_bresp   ,
    output          o_bvalid  ,
    input           i_bready  ,
    input  [3:0]    i_arid    ,
    input  [31:0]   i_araddr  ,
    input  [3:0]    i_arlen   ,
    input  [2:0]    i_arsize  ,
    input  [1:0]    i_arburst ,
    input  [1:0]    i_arlock  ,
    input  [3:0]    i_arcache ,
    input  [2:0]    i_arprot  ,
    input           i_arvalid ,
    output          o_arready ,
    output [3:0]    o_rid     ,
    output [127:0]  o_rdata   ,
    output [1:0]    o_rresp   ,
    output          o_rlast   ,
    output          o_rvalid  ,
    input           i_rready  ,

    output          o_cs      ,
    output [31:0]   o_addr    ,
    output [31:0]   o_data    ,
    input  [31:0]   i_data
);


endmodule