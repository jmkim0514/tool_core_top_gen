//==============================================================================
//
// Project : MVP
//
// Verilog RTL(Behavioral) model
//
// This confidential and proprietary source code may be used only as authorized
// by a licensing agreement from ALPHAHOLDINGS Limited. The entire notice above
// must be reproduced on all authorized copies and copies may only be made to
// the extent permitted by a licensing agreement from ALPHAHOLDINGS Limited.
//
// COPYRIGHT (C) ALPHAHOLDINGS, inc. 2022
//
//==============================================================================
// File name : ddr_hpdf
// Version : v1.1
// Description :
// Simulator : NC Verilog
// Created by : yhsim
// Date : 2023-11-03  15:16
//==============================================================================

module ddr_hpdf (
    input              i_test_bypass,
    input              i_rstn_peri2ddr,
    input              i_clk_peri2ddr,
    input              i_clk_xtal_y,
    input              i_clk_main2ddr,
    input              i_scan_clk,
    input              i_scan_mode,
    input              i_test_rstn,
    input   [  1:  0]  i_pll2651_mode,
    input   [  5:  0]  t_ddr_pll_p,
    input   [  8:  0]  t_ddr_pll_m,
    input   [  2:  0]  t_ddr_pll_s,
    input   [ 15:  0]  t_ddr_pll_k,
    input   [  4:  0]  t_ddr_pll_extafc,
    input   [  7:  0]  t_ddr_pll_mfr,
    input   [  5:  0]  t_ddr_pll_mrr,
    input   [  1:  0]  t_ddr_pll_sel_pf,
    input   [  1:  0]  t_ddr_pll_icp,
    input              t_ddr_pll_pbias_ctrl,
    input              t_ddr_pll_pbias_ctrl_en,
    input              t_ddr_pll_vco_boost,
    input              t_ddr_pll_resetb,
    input              t_ddr_pll_fsel,
    input              t_ddr_pll_fvco_en,
    input              t_ddr_pll_bypass,
    input              t_ddr_pll_sscg_en,
    input              t_ddr_pll_afc_enb,
    input              t_ddr_pll_afcinit_sel,
    input              t_ddr_pll_fout_mask,
    input              t_ddr_pll_lrd_en,
    input   [  5:  0]  sr_ddr_pll_p,
    input   [  8:  0]  sr_ddr_pll_m,
    input   [  2:  0]  sr_ddr_pll_s,
    input   [ 15:  0]  sr_ddr_pll_k,
    output             t_ddr_pll_fout,
    output             t_ddr_pll_fvco_out,
    output  [  4:  0]  t_ddr_pll_afc_code,
    input   [  8:  0]  i_awid_main2ddr_s1,
    input   [ 31:  0]  i_awaddr_main2ddr_s1,
    input   [  7:  0]  i_awlen_main2ddr_s1,
    input   [  2:  0]  i_awsize_main2ddr_s1,
    input   [  1:  0]  i_awburst_main2ddr_s1,
    input              i_awlock_main2ddr_s1,
    input   [  3:  0]  i_awcache_main2ddr_s1,
    input   [  2:  0]  i_awprot_main2ddr_s1,
    input              i_awvalid_main2ddr_s1,
    output             o_awready_main2ddr_s1,
    input   [127:  0]  i_wdata_main2ddr_s1,
    input   [ 15:  0]  i_wstrb_main2ddr_s1,
    input              i_wlast_main2ddr_s1,
    input              i_wvalid_main2ddr_s1,
    output             o_wready_main2ddr_s1,
    output  [  8:  0]  o_bid_main2ddr_s1,
    output  [  1:  0]  o_bresp_main2ddr_s1,
    output             o_bvalid_main2ddr_s1,
    input              i_bready_main2ddr_s1,
    input   [  8:  0]  i_arid_main2ddr_s1,
    input   [ 31:  0]  i_araddr_main2ddr_s1,
    input   [  7:  0]  i_arlen_main2ddr_s1,
    input   [  2:  0]  i_arsize_main2ddr_s1,
    input   [  1:  0]  i_arburst_main2ddr_s1,
    input              i_arlock_main2ddr_s1,
    input   [  3:  0]  i_arcache_main2ddr_s1,
    input   [  2:  0]  i_arprot_main2ddr_s1,
    input              i_arvalid_main2ddr_s1,
    output             o_arready_main2ddr_s1,
    output  [  8:  0]  o_rid_main2ddr_s1,
    output  [127:  0]  o_rdata_main2ddr_s1,
    output  [  1:  0]  o_rresp_main2ddr_s1,
    output             o_rlast_main2ddr_s1,
    output             o_rvalid_main2ddr_s1,
    input              i_rready_main2ddr_s1,
    input   [  8:  0]  i_awid_main2ddr_s2,
    input   [ 31:  0]  i_awaddr_main2ddr_s2,
    input   [  7:  0]  i_awlen_main2ddr_s2,
    input   [  2:  0]  i_awsize_main2ddr_s2,
    input   [  1:  0]  i_awburst_main2ddr_s2,
    input              i_awlock_main2ddr_s2,
    input   [  3:  0]  i_awcache_main2ddr_s2,
    input   [  2:  0]  i_awprot_main2ddr_s2,
    input              i_awvalid_main2ddr_s2,
    output             o_awready_main2ddr_s2,
    input   [127:  0]  i_wdata_main2ddr_s2,
    input   [ 15:  0]  i_wstrb_main2ddr_s2,
    input              i_wlast_main2ddr_s2,
    input              i_wvalid_main2ddr_s2,
    output             o_wready_main2ddr_s2,
    output  [  8:  0]  o_bid_main2ddr_s2,
    output  [  1:  0]  o_bresp_main2ddr_s2,
    output             o_bvalid_main2ddr_s2,
    input              i_bready_main2ddr_s2,
    input   [  8:  0]  i_arid_main2ddr_s2,
    input   [ 31:  0]  i_araddr_main2ddr_s2,
    input   [  7:  0]  i_arlen_main2ddr_s2,
    input   [  2:  0]  i_arsize_main2ddr_s2,
    input   [  1:  0]  i_arburst_main2ddr_s2,
    input              i_arlock_main2ddr_s2,
    input   [  3:  0]  i_arcache_main2ddr_s2,
    input   [  2:  0]  i_arprot_main2ddr_s2,
    input              i_arvalid_main2ddr_s2,
    output             o_arready_main2ddr_s2,
    output  [  8:  0]  o_rid_main2ddr_s2,
    output  [127:  0]  o_rdata_main2ddr_s2,
    output  [  1:  0]  o_rresp_main2ddr_s2,
    output             o_rlast_main2ddr_s2,
    output             o_rvalid_main2ddr_s2,
    input              i_rready_main2ddr_s2,
    input   [  8:  0]  i_awid_main2ddr_s3,
    input   [ 31:  0]  i_awaddr_main2ddr_s3,
    input   [  7:  0]  i_awlen_main2ddr_s3,
    input   [  2:  0]  i_awsize_main2ddr_s3,
    input   [  1:  0]  i_awburst_main2ddr_s3,
    input              i_awlock_main2ddr_s3,
    input   [  3:  0]  i_awcache_main2ddr_s3,
    input   [  2:  0]  i_awprot_main2ddr_s3,
    input              i_awvalid_main2ddr_s3,
    output             o_awready_main2ddr_s3,
    input   [127:  0]  i_wdata_main2ddr_s3,
    input   [ 15:  0]  i_wstrb_main2ddr_s3,
    input              i_wlast_main2ddr_s3,
    input              i_wvalid_main2ddr_s3,
    output             o_wready_main2ddr_s3,
    output  [  8:  0]  o_bid_main2ddr_s3,
    output  [  1:  0]  o_bresp_main2ddr_s3,
    output             o_bvalid_main2ddr_s3,
    input              i_bready_main2ddr_s3,
    input   [  8:  0]  i_arid_main2ddr_s3,
    input   [ 31:  0]  i_araddr_main2ddr_s3,
    input   [  7:  0]  i_arlen_main2ddr_s3,
    input   [  2:  0]  i_arsize_main2ddr_s3,
    input   [  1:  0]  i_arburst_main2ddr_s3,
    input              i_arlock_main2ddr_s3,
    input   [  3:  0]  i_arcache_main2ddr_s3,
    input   [  2:  0]  i_arprot_main2ddr_s3,
    input              i_arvalid_main2ddr_s3,
    output             o_arready_main2ddr_s3,
    output  [  8:  0]  o_rid_main2ddr_s3,
    output  [127:  0]  o_rdata_main2ddr_s3,
    output  [  1:  0]  o_rresp_main2ddr_s3,
    output             o_rlast_main2ddr_s3,
    output             o_rvalid_main2ddr_s3,
    input              i_rready_main2ddr_s3,
    output             o_irq_asp,
    output             o_irq_overtemp,
    output             o_irq_hightemp,
    output             o_irq_cooldown,
    inout              DDR_VREF0,
    inout              DDR_VREF1,
    input              DDR_MEM_CKEIN,
    output             DDR_MEM_CK_P,
    output             DDR_MEM_CK_N,
    inout   [  1:  0]  DDR_MEM_CKE,
    inout              DDR_MEM_RESET_N,
    inout   [  1:  0]  DDR_MEM_ODT,
    inout   [  1:  0]  DDR_MEM_CSN,
    inout              DDR_MEM_RASN,
    inout              DDR_MEM_CASN,
    inout              DDR_MEM_WEN,
    inout   [  2:  0]  DDR_MEM_BA,
    inout   [ 15:  0]  DDR_MEM_A,
    inout   [ 31:  0]  DDR_MEM_DQ,
    inout   [  3:  0]  DDR_MEM_DM,
    inout   [  3:  0]  DDR_MEM_DQS_P,
    inout   [  3:  0]  DDR_MEM_DQS_N,
    inout              DDR_ZQ,
    input              t_ddr_phy_phy_y,
    input              t_ddr_phy_scan_y,
    input              t_ddr_phy_nand_y,
    input   [  2:  0]  t_ddr_phy_run_y,
    input              t_ddr_phy_mux_y,
    input              t_ddr_phy_highz_y,
    input              t_ddr_phy_ext_en_y,
    input              t_ddr_phy_ext_out_y,
    input              t_ddr_phy_ext_read_y,
    input              t_ddr_phy_ext_cmosrcv_y,
    input              t_ddr_phy_ext_zq_force_y,
    input   [  2:  0]  t_ddr_phy_ext_zq_force_impp_y,
    input   [  2:  0]  t_ddr_phy_ext_zq_force_impn_y,
    input   [  2:  0]  t_ddr_phy_ext_zq_mode_dds_y,
    input              t_ddr_phy_ext_dfdqs_y,
    input   [  3:  0]  t_ddr_phy_ext_ref_y,
    input   [  7:  0]  t_ddr_phy_ext_offsetc_y,
    input              t_ddr_phy_ext_rdlvl_en_y,
    input              t_ddr_phy_ext_rdlvl_wr_en_y,
    input              t_ddr_phy_ext_gatelvl_en_y,
    input              t_ddr_phy_ext_write_lvl_en_y,
    input              t_ddr_phy_ext_ca_cal_en_y,
    input   [  3:  0]  t_ddr_phy_ext_mode_y,
    input   [  4:  0]  t_ddr_phy_start_y,
    input   [  3:  0]  t_ddr_phy_ext_rdlvl_incr_adj_y,
    output             t_ddr_phy_ctrl_div_out_400_a,
    output             t_ddr_phy_ctrl_div_out_800_a,
    output             t_ddr_phy_ext_zq_end_a,
    output  [  8:  0]  t_ddr_phy_ext_lock_value_a,
    output             t_ddr_phy_ext_clock_a,
    output             t_ddr_phy_ext_flock_a,
    output             t_ddr_phy_ext_locked_a,
    output             t_ddr_phy_ext_init_complete_a,
    output  [  3:  0]  t_ddr_phy_ext_rdlvl_vwmc_a,
    output  [  4:  0]  t_ddr_phy_err_a,
    output  [  4:  0]  t_ddr_phy_oky_a,
    input              test_se,
    input   [ 35:  0]  test_si,
    output  [ 35:  0]  test_so,
    input              i_psel_ddr_m0_deco,
    input              i_penable_ddr_m0_deco,
    input   [ 31:  0]  i_paddr_ddr_m0_deco,
    input              i_pwrite_ddr_m0_deco,
    input   [ 31:  0]  i_pwdata_ddr_m0_deco,
    output  [ 31:  0]  o_prdata_ddr_m0_deco,
    output             o_pready_ddr_m0_deco,
    output             o_pslverr_ddr_m0_deco
);

    wire             ddr_crm_o_pll_resetb;
    wire             ddr_crm_o_pll_bypass;
    wire    [  5:0]  ddr_crm_o_pll_p;
    wire    [  8:0]  ddr_crm_o_pll_m;
    wire    [  2:0]  ddr_crm_o_pll_s;
    wire    [ 15:0]  ddr_crm_o_pll_k;
    wire    [  4:0]  ddr_crm_o_pll_extafc;
    wire    [  7:0]  ddr_crm_o_pll_mfr;
    wire    [  5:0]  ddr_crm_o_pll_mrr;
    wire    [  1:0]  ddr_crm_o_pll_sel_pf;
    wire    [  1:0]  ddr_crm_o_pll_icp;
    wire             ddr_crm_o_pll_pbias_ctrl;
    wire             ddr_crm_o_pll_pbias_ctrl_en;
    wire             ddr_crm_o_pll_vco_boost;
    wire             ddr_crm_o_pll_fsel;
    wire             ddr_crm_o_pll_fvco_en;
    wire             ddr_crm_o_pll_sscg_en;
    wire             ddr_crm_o_pll_afc_enb;
    wire             ddr_crm_o_pll_afcinit_sel;
    wire             ddr_crm_o_pll_fout_mask;
    wire             ddr_crm_o_pll_lrd_en;
    wire             ddr_crm_o_clk_ddr_ref;
    wire             ddr_crm_o_rstn_ddr_ref;
    wire             ddr_crm_o_clk_peri2ddr;
    wire             ddr_crm_o_rstn_peri2ddr;
    wire             ddr_crm_o_sclk_omc;
    wire             ddr_crm_o_srstn_omc;
    wire             ddr_crm_o_sclk_ddr_phy;
    wire             ddr_crm_o_srstn_ddr_phy;
    wire             ddr_crm_o_mclk_ddr_phy;
    wire             ddr_crm_o_mrstn_ddr_phy;
    wire             ddr_crm_o_clk_ddr_phym;
    wire             ddr_crm_o_mclk_omc;
    wire             ddr_crm_o_mrstn_omc;
    wire             ddr_crm_o_clk_main2ddr;
    wire             ddr_crm_o_rstn_main2ddr;
    wire             pll_top_ddr_o_fout;
    wire             pll_top_ddr_o_fvco_out;
    wire    [  4:0]  pll_top_ddr_o_afc_code;
    wire    [ 10:0]  ddr_bus_awid_ddr_m0;
    wire    [ 31:0]  ddr_bus_awaddr_ddr_m0;
    wire    [  7:0]  ddr_bus_awlen_ddr_m0;
    wire    [  2:0]  ddr_bus_awsize_ddr_m0;
    wire    [  1:0]  ddr_bus_awburst_ddr_m0;
    wire             ddr_bus_awlock_ddr_m0;
    wire    [  3:0]  ddr_bus_awcache_ddr_m0;
    wire    [  2:0]  ddr_bus_awprot_ddr_m0;
    wire             ddr_bus_awvalid_ddr_m0;
    wire             ddr_bus_awready_ddr_m0;
    wire    [127:0]  ddr_bus_wdata_ddr_m0;
    wire    [ 15:0]  ddr_bus_wstrb_ddr_m0;
    wire             ddr_bus_wlast_ddr_m0;
    wire             ddr_bus_wvalid_ddr_m0;
    wire             ddr_bus_wready_ddr_m0;
    wire    [ 10:0]  ddr_bus_bid_ddr_m0;
    wire    [  1:0]  ddr_bus_bresp_ddr_m0;
    wire             ddr_bus_bvalid_ddr_m0;
    wire             ddr_bus_bready_ddr_m0;
    wire    [ 10:0]  ddr_bus_arid_ddr_m0;
    wire    [ 31:0]  ddr_bus_araddr_ddr_m0;
    wire    [  7:0]  ddr_bus_arlen_ddr_m0;
    wire    [  2:0]  ddr_bus_arsize_ddr_m0;
    wire    [  1:0]  ddr_bus_arburst_ddr_m0;
    wire             ddr_bus_arlock_ddr_m0;
    wire    [  3:0]  ddr_bus_arcache_ddr_m0;
    wire    [  2:0]  ddr_bus_arprot_ddr_m0;
    wire             ddr_bus_arvalid_ddr_m0;
    wire             ddr_bus_arready_ddr_m0;
    wire    [ 10:0]  ddr_bus_rid_ddr_m0;
    wire    [127:0]  ddr_bus_rdata_ddr_m0;
    wire    [  1:0]  ddr_bus_rresp_ddr_m0;
    wire             ddr_bus_rlast_ddr_m0;
    wire             ddr_bus_rvalid_ddr_m0;
    wire             ddr_bus_rready_ddr_m0;
    wire             ddr_sub_o_clk_dfi;
    wire             ddr_sub_o_psel_ddr_crm;
    wire             ddr_sub_o_penable_ddr_crm;
    wire    [ 11:0]  ddr_sub_o_paddr_ddr_crm;
    wire             ddr_sub_o_pwrite_ddr_crm;
    wire    [ 31:0]  ddr_sub_o_pwdata_ddr_crm;
    wire    [ 31:0]  ddr_sub_i_prdata_ddr_crm;
    wire    [ 31:0]  ddr_sub_o_haddr_ddr_bus_gpv;
    wire    [  2:0]  ddr_sub_o_hburst_ddr_bus_gpv;
    wire    [  2:0]  ddr_sub_o_hsize_ddr_bus_gpv;
    wire    [  1:0]  ddr_sub_o_htrans_ddr_bus_gpv;
    wire    [ 31:0]  ddr_sub_o_hwdata_ddr_bus_gpv;
    wire             ddr_sub_o_hwrite_ddr_bus_gpv;
    wire    [ 31:0]  ddr_sub_i_hrdata_ddr_bus_gpv;
    wire             ddr_sub_i_hreadyout_ddr_bus_gpv;
    wire             ddr_sub_i_hresp_ddr_bus_gpv;

    assign  t_ddr_pll_afc_code[4:0] = pll_top_ddr_o_afc_code[4:0];
    assign  t_ddr_pll_fout = pll_top_ddr_o_fout;
    assign  t_ddr_pll_fvco_out = pll_top_ddr_o_fvco_out;

    mvp_crm_ddr u_ddr_crm (
        .i_test_bypass                 (i_test_bypass),
        .i_rstn_peri                   (i_rstn_peri2ddr),
        .i_apb_pclk                    (i_clk_peri2ddr),
        .i_apb_prstn                   (i_rstn_peri2ddr),
        .i_apb_psel                    (ddr_sub_o_psel_ddr_crm),
        .i_apb_penable                 (ddr_sub_o_penable_ddr_crm),
        .i_apb_pwrite                  (ddr_sub_o_pwrite_ddr_crm),
        .i_apb_paddr                   (ddr_sub_o_paddr_ddr_crm),
        .i_apb_pwdata                  (ddr_sub_o_pwdata_ddr_crm),
        .o_apb_prdata                  (ddr_sub_i_prdata_ddr_crm),
        .o_pll_resetb                  (ddr_crm_o_pll_resetb),
        .o_pll_bypass                  (ddr_crm_o_pll_bypass),
        .o_pll_p                       (ddr_crm_o_pll_p),
        .o_pll_m                       (ddr_crm_o_pll_m),
        .o_pll_s                       (ddr_crm_o_pll_s),
        .o_pll_k                       (ddr_crm_o_pll_k),
        .o_pll_extafc                  (ddr_crm_o_pll_extafc),
        .o_pll_mfr                     (ddr_crm_o_pll_mfr),
        .o_pll_mrr                     (ddr_crm_o_pll_mrr),
        .o_pll_sel_pf                  (ddr_crm_o_pll_sel_pf),
        .o_pll_icp                     (ddr_crm_o_pll_icp),
        .o_pll_pbias_ctrl              (ddr_crm_o_pll_pbias_ctrl),
        .o_pll_pbias_ctrl_en           (ddr_crm_o_pll_pbias_ctrl_en),
        .o_pll_vco_boost               (ddr_crm_o_pll_vco_boost),
        .o_pll_fsel                    (ddr_crm_o_pll_fsel),
        .o_pll_fvco_en                 (ddr_crm_o_pll_fvco_en),
        .o_pll_sscg_en                 (ddr_crm_o_pll_sscg_en),
        .o_pll_afc_enb                 (ddr_crm_o_pll_afc_enb),
        .o_pll_afcinit_sel             (ddr_crm_o_pll_afcinit_sel),
        .o_pll_fout_mask               (ddr_crm_o_pll_fout_mask),
        .o_pll_lrd_en                  (ddr_crm_o_pll_lrd_en),
        .i_pll_fvco_out                (pll_top_ddr_o_fvco_out),
        .i_pll_afc_code                (pll_top_ddr_o_afc_code),
        .i_clk_xtal_y                  (i_clk_xtal_y),
        .i_clk_peri2ddr                (i_clk_peri2ddr),
        .i_clk_pll_ddr                 (pll_top_ddr_o_fout),
        .i_clk_dfi_phy                 (ddr_sub_o_clk_dfi),
        .i_clk_main2ddr                (i_clk_main2ddr),
        .o_clk_ddr_ref                 (ddr_crm_o_clk_ddr_ref),
        .o_rstn_ddr_ref                (ddr_crm_o_rstn_ddr_ref),
        .o_clk_peri2ddr                (ddr_crm_o_clk_peri2ddr),
        .o_rstn_peri2ddr               (ddr_crm_o_rstn_peri2ddr),
        .o_sclk_omc                    (ddr_crm_o_sclk_omc),
        .o_srstn_omc                   (ddr_crm_o_srstn_omc),
        .o_sclk_ddr_phy                (ddr_crm_o_sclk_ddr_phy),
        .o_srstn_ddr_phy               (ddr_crm_o_srstn_ddr_phy),
        .o_mclk_ddr_phy                (ddr_crm_o_mclk_ddr_phy),
        .o_mrstn_ddr_phy               (ddr_crm_o_mrstn_ddr_phy),
        .o_clk_ddr_phym                (ddr_crm_o_clk_ddr_phym),
        .o_mclk_omc                    (ddr_crm_o_mclk_omc),
        .o_mrstn_omc                   (ddr_crm_o_mrstn_omc),
        .o_clk_main2ddr                (ddr_crm_o_clk_main2ddr),
        .o_rstn_main2ddr               (ddr_crm_o_rstn_main2ddr),
        .i_scan_clk                    (i_scan_clk),
        .i_scan_mode                   (i_scan_mode),
        .i_scan_rstn                   (i_test_rstn)
    );

    tmux_sf_pll2651x_ln28lpp_5000 u_pll_top_ddr (
        .i_tmode                       (i_pll2651_mode),
        .i_norm_p                      (ddr_crm_o_pll_p),
        .i_norm_m                      (ddr_crm_o_pll_m),
        .i_norm_s                      (ddr_crm_o_pll_s),
        .i_norm_k                      (ddr_crm_o_pll_k),
        .i_norm_extafc                 (ddr_crm_o_pll_extafc),
        .i_norm_mfr                    (ddr_crm_o_pll_mfr),
        .i_norm_mrr                    (ddr_crm_o_pll_mrr),
        .i_norm_sel_pf                 (ddr_crm_o_pll_sel_pf),
        .i_norm_icp                    (ddr_crm_o_pll_icp),
        .i_norm_pbias_ctrl             (ddr_crm_o_pll_pbias_ctrl),
        .i_norm_pbias_ctrl_en          (ddr_crm_o_pll_pbias_ctrl_en),
        .i_norm_vco_boost              (ddr_crm_o_pll_vco_boost),
        .i_norm_fin                    (i_clk_xtal_y),
        .i_norm_resetb                 (ddr_crm_o_pll_resetb),
        .i_norm_fsel                   (ddr_crm_o_pll_fsel),
        .i_norm_fvco_en                (ddr_crm_o_pll_fvco_en),
        .i_norm_bypass                 (ddr_crm_o_pll_bypass),
        .i_norm_sscg_en                (ddr_crm_o_pll_sscg_en),
        .i_norm_afc_enb                (ddr_crm_o_pll_afc_enb),
        .i_norm_afcinit_sel            (ddr_crm_o_pll_afcinit_sel),
        .i_norm_fout_mask              (ddr_crm_o_pll_fout_mask),
        .i_norm_lrd_en                 (ddr_crm_o_pll_lrd_en),
        .i_test0_p                     (t_ddr_pll_p),
        .i_test0_m                     (t_ddr_pll_m),
        .i_test0_s                     (t_ddr_pll_s),
        .i_test0_k                     (t_ddr_pll_k),
        .i_test0_extafc                (t_ddr_pll_extafc),
        .i_test0_mfr                   (t_ddr_pll_mfr),
        .i_test0_mrr                   (t_ddr_pll_mrr),
        .i_test0_sel_pf                (t_ddr_pll_sel_pf),
        .i_test0_icp                   (t_ddr_pll_icp),
        .i_test0_pbias_ctrl            (t_ddr_pll_pbias_ctrl),
        .i_test0_pbias_ctrl_en         (t_ddr_pll_pbias_ctrl_en),
        .i_test0_vco_boost             (t_ddr_pll_vco_boost),
        .i_test0_fin                   (i_clk_xtal_y),
        .i_test0_resetb                (t_ddr_pll_resetb),
        .i_test0_fsel                  (t_ddr_pll_fsel),
        .i_test0_fvco_en               (t_ddr_pll_fvco_en),
        .i_test0_bypass                (t_ddr_pll_bypass),
        .i_test0_sscg_en               (t_ddr_pll_sscg_en),
        .i_test0_afc_enb               (t_ddr_pll_afc_enb),
        .i_test0_afcinit_sel           (t_ddr_pll_afcinit_sel),
        .i_test0_fout_mask             (t_ddr_pll_fout_mask),
        .i_test0_lrd_en                (t_ddr_pll_lrd_en),
        .i_test1_p                     (sr_ddr_pll_p),
        .i_test1_m                     (sr_ddr_pll_m),
        .i_test1_s                     (sr_ddr_pll_s),
        .i_test1_k                     (sr_ddr_pll_k),
        .i_test1_extafc                (5'h0),
        .i_test1_mfr                   (8'h8),
        .i_test1_mrr                   (6'h30),
        .i_test1_sel_pf                (2'h0),
        .i_test1_icp                   (2'h0),
        .i_test1_pbias_ctrl            (1'h0),
        .i_test1_pbias_ctrl_en         (1'h0),
        .i_test1_vco_boost             (1'h1),
        .i_test1_fin                   (i_clk_xtal_y),
        .i_test1_resetb                (t_ddr_pll_resetb),
        .i_test1_fsel                  (1'h0),
        .i_test1_fvco_en               (1'h0),
        .i_test1_bypass                (1'h0),
        .i_test1_sscg_en               (1'h0),
        .i_test1_afc_enb               (1'h0),
        .i_test1_afcinit_sel           (1'h1),
        .i_test1_fout_mask             (1'h0),
        .i_test1_lrd_en                (1'h0),
        .o_fout                        (pll_top_ddr_o_fout),
        .o_fvco_out                    (pll_top_ddr_o_fvco_out),
        .o_afc_code                    (pll_top_ddr_o_afc_code)
    );

    nic400_ddr_bus_r0p00 u_ddr_bus (
        .awid_ddr_m0                   (ddr_bus_awid_ddr_m0),
        .awaddr_ddr_m0                 (ddr_bus_awaddr_ddr_m0),
        .awlen_ddr_m0                  (ddr_bus_awlen_ddr_m0),
        .awsize_ddr_m0                 (ddr_bus_awsize_ddr_m0),
        .awburst_ddr_m0                (ddr_bus_awburst_ddr_m0),
        .awlock_ddr_m0                 (ddr_bus_awlock_ddr_m0),
        .awcache_ddr_m0                (ddr_bus_awcache_ddr_m0),
        .awprot_ddr_m0                 (ddr_bus_awprot_ddr_m0),
        .awvalid_ddr_m0                (ddr_bus_awvalid_ddr_m0),
        .awready_ddr_m0                (ddr_bus_awready_ddr_m0),
        .wdata_ddr_m0                  (ddr_bus_wdata_ddr_m0),
        .wstrb_ddr_m0                  (ddr_bus_wstrb_ddr_m0),
        .wlast_ddr_m0                  (ddr_bus_wlast_ddr_m0),
        .wvalid_ddr_m0                 (ddr_bus_wvalid_ddr_m0),
        .wready_ddr_m0                 (ddr_bus_wready_ddr_m0),
        .bid_ddr_m0                    (ddr_bus_bid_ddr_m0),
        .bresp_ddr_m0                  (ddr_bus_bresp_ddr_m0),
        .bvalid_ddr_m0                 (ddr_bus_bvalid_ddr_m0),
        .bready_ddr_m0                 (ddr_bus_bready_ddr_m0),
        .arid_ddr_m0                   (ddr_bus_arid_ddr_m0),
        .araddr_ddr_m0                 (ddr_bus_araddr_ddr_m0),
        .arlen_ddr_m0                  (ddr_bus_arlen_ddr_m0),
        .arsize_ddr_m0                 (ddr_bus_arsize_ddr_m0),
        .arburst_ddr_m0                (ddr_bus_arburst_ddr_m0),
        .arlock_ddr_m0                 (ddr_bus_arlock_ddr_m0),
        .arcache_ddr_m0                (ddr_bus_arcache_ddr_m0),
        .arprot_ddr_m0                 (ddr_bus_arprot_ddr_m0),
        .arvalid_ddr_m0                (ddr_bus_arvalid_ddr_m0),
        .arready_ddr_m0                (ddr_bus_arready_ddr_m0),
        .rid_ddr_m0                    (ddr_bus_rid_ddr_m0),
        .rdata_ddr_m0                  (ddr_bus_rdata_ddr_m0),
        .rresp_ddr_m0                  (ddr_bus_rresp_ddr_m0),
        .rlast_ddr_m0                  (ddr_bus_rlast_ddr_m0),
        .rvalid_ddr_m0                 (ddr_bus_rvalid_ddr_m0),
        .rready_ddr_m0                 (ddr_bus_rready_ddr_m0),
        .awid_main2ddr_s1              (i_awid_main2ddr_s1),
        .awaddr_main2ddr_s1            (i_awaddr_main2ddr_s1),
        .awlen_main2ddr_s1             (i_awlen_main2ddr_s1),
        .awsize_main2ddr_s1            (i_awsize_main2ddr_s1),
        .awburst_main2ddr_s1           (i_awburst_main2ddr_s1),
        .awlock_main2ddr_s1            (i_awlock_main2ddr_s1),
        .awcache_main2ddr_s1           (i_awcache_main2ddr_s1),
        .awprot_main2ddr_s1            (i_awprot_main2ddr_s1),
        .awvalid_main2ddr_s1           (i_awvalid_main2ddr_s1),
        .awready_main2ddr_s1           (o_awready_main2ddr_s1),
        .wdata_main2ddr_s1             (i_wdata_main2ddr_s1),
        .wstrb_main2ddr_s1             (i_wstrb_main2ddr_s1),
        .wlast_main2ddr_s1             (i_wlast_main2ddr_s1),
        .wvalid_main2ddr_s1            (i_wvalid_main2ddr_s1),
        .wready_main2ddr_s1            (o_wready_main2ddr_s1),
        .bid_main2ddr_s1               (o_bid_main2ddr_s1),
        .bresp_main2ddr_s1             (o_bresp_main2ddr_s1),
        .bvalid_main2ddr_s1            (o_bvalid_main2ddr_s1),
        .bready_main2ddr_s1            (i_bready_main2ddr_s1),
        .arid_main2ddr_s1              (i_arid_main2ddr_s1),
        .araddr_main2ddr_s1            (i_araddr_main2ddr_s1),
        .arlen_main2ddr_s1             (i_arlen_main2ddr_s1),
        .arsize_main2ddr_s1            (i_arsize_main2ddr_s1),
        .arburst_main2ddr_s1           (i_arburst_main2ddr_s1),
        .arlock_main2ddr_s1            (i_arlock_main2ddr_s1),
        .arcache_main2ddr_s1           (i_arcache_main2ddr_s1),
        .arprot_main2ddr_s1            (i_arprot_main2ddr_s1),
        .arvalid_main2ddr_s1           (i_arvalid_main2ddr_s1),
        .arready_main2ddr_s1           (o_arready_main2ddr_s1),
        .rid_main2ddr_s1               (o_rid_main2ddr_s1),
        .rdata_main2ddr_s1             (o_rdata_main2ddr_s1),
        .rresp_main2ddr_s1             (o_rresp_main2ddr_s1),
        .rlast_main2ddr_s1             (o_rlast_main2ddr_s1),
        .rvalid_main2ddr_s1            (o_rvalid_main2ddr_s1),
        .rready_main2ddr_s1            (i_rready_main2ddr_s1),
        .awid_main2ddr_s2              (i_awid_main2ddr_s2),
        .awaddr_main2ddr_s2            (i_awaddr_main2ddr_s2),
        .awlen_main2ddr_s2             (i_awlen_main2ddr_s2),
        .awsize_main2ddr_s2            (i_awsize_main2ddr_s2),
        .awburst_main2ddr_s2           (i_awburst_main2ddr_s2),
        .awlock_main2ddr_s2            (i_awlock_main2ddr_s2),
        .awcache_main2ddr_s2           (i_awcache_main2ddr_s2),
        .awprot_main2ddr_s2            (i_awprot_main2ddr_s2),
        .awvalid_main2ddr_s2           (i_awvalid_main2ddr_s2),
        .awready_main2ddr_s2           (o_awready_main2ddr_s2),
        .wdata_main2ddr_s2             (i_wdata_main2ddr_s2),
        .wstrb_main2ddr_s2             (i_wstrb_main2ddr_s2),
        .wlast_main2ddr_s2             (i_wlast_main2ddr_s2),
        .wvalid_main2ddr_s2            (i_wvalid_main2ddr_s2),
        .wready_main2ddr_s2            (o_wready_main2ddr_s2),
        .bid_main2ddr_s2               (o_bid_main2ddr_s2),
        .bresp_main2ddr_s2             (o_bresp_main2ddr_s2),
        .bvalid_main2ddr_s2            (o_bvalid_main2ddr_s2),
        .bready_main2ddr_s2            (i_bready_main2ddr_s2),
        .arid_main2ddr_s2              (i_arid_main2ddr_s2),
        .araddr_main2ddr_s2            (i_araddr_main2ddr_s2),
        .arlen_main2ddr_s2             (i_arlen_main2ddr_s2),
        .arsize_main2ddr_s2            (i_arsize_main2ddr_s2),
        .arburst_main2ddr_s2           (i_arburst_main2ddr_s2),
        .arlock_main2ddr_s2            (i_arlock_main2ddr_s2),
        .arcache_main2ddr_s2           (i_arcache_main2ddr_s2),
        .arprot_main2ddr_s2            (i_arprot_main2ddr_s2),
        .arvalid_main2ddr_s2           (i_arvalid_main2ddr_s2),
        .arready_main2ddr_s2           (o_arready_main2ddr_s2),
        .rid_main2ddr_s2               (o_rid_main2ddr_s2),
        .rdata_main2ddr_s2             (o_rdata_main2ddr_s2),
        .rresp_main2ddr_s2             (o_rresp_main2ddr_s2),
        .rlast_main2ddr_s2             (o_rlast_main2ddr_s2),
        .rvalid_main2ddr_s2            (o_rvalid_main2ddr_s2),
        .rready_main2ddr_s2            (i_rready_main2ddr_s2),
        .awid_main2ddr_s3              (i_awid_main2ddr_s3),
        .awaddr_main2ddr_s3            (i_awaddr_main2ddr_s3),
        .awlen_main2ddr_s3             (i_awlen_main2ddr_s3),
        .awsize_main2ddr_s3            (i_awsize_main2ddr_s3),
        .awburst_main2ddr_s3           (i_awburst_main2ddr_s3),
        .awlock_main2ddr_s3            (i_awlock_main2ddr_s3),
        .awcache_main2ddr_s3           (i_awcache_main2ddr_s3),
        .awprot_main2ddr_s3            (i_awprot_main2ddr_s3),
        .awvalid_main2ddr_s3           (i_awvalid_main2ddr_s3),
        .awready_main2ddr_s3           (o_awready_main2ddr_s3),
        .wdata_main2ddr_s3             (i_wdata_main2ddr_s3),
        .wstrb_main2ddr_s3             (i_wstrb_main2ddr_s3),
        .wlast_main2ddr_s3             (i_wlast_main2ddr_s3),
        .wvalid_main2ddr_s3            (i_wvalid_main2ddr_s3),
        .wready_main2ddr_s3            (o_wready_main2ddr_s3),
        .bid_main2ddr_s3               (o_bid_main2ddr_s3),
        .bresp_main2ddr_s3             (o_bresp_main2ddr_s3),
        .bvalid_main2ddr_s3            (o_bvalid_main2ddr_s3),
        .bready_main2ddr_s3            (i_bready_main2ddr_s3),
        .arid_main2ddr_s3              (i_arid_main2ddr_s3),
        .araddr_main2ddr_s3            (i_araddr_main2ddr_s3),
        .arlen_main2ddr_s3             (i_arlen_main2ddr_s3),
        .arsize_main2ddr_s3            (i_arsize_main2ddr_s3),
        .arburst_main2ddr_s3           (i_arburst_main2ddr_s3),
        .arlock_main2ddr_s3            (i_arlock_main2ddr_s3),
        .arcache_main2ddr_s3           (i_arcache_main2ddr_s3),
        .arprot_main2ddr_s3            (i_arprot_main2ddr_s3),
        .arvalid_main2ddr_s3           (i_arvalid_main2ddr_s3),
        .arready_main2ddr_s3           (o_arready_main2ddr_s3),
        .rid_main2ddr_s3               (o_rid_main2ddr_s3),
        .rdata_main2ddr_s3             (o_rdata_main2ddr_s3),
        .rresp_main2ddr_s3             (o_rresp_main2ddr_s3),
        .rlast_main2ddr_s3             (o_rlast_main2ddr_s3),
        .rvalid_main2ddr_s3            (o_rvalid_main2ddr_s3),
        .rready_main2ddr_s3            (i_rready_main2ddr_s3),
        .haddr_ddr_bus_gpv_s0          (ddr_sub_o_haddr_ddr_bus_gpv),
        .hburst_ddr_bus_gpv_s0         (ddr_sub_o_hburst_ddr_bus_gpv),
        .hprot_ddr_bus_gpv_s0          (4'h0),
        .hsize_ddr_bus_gpv_s0          (ddr_sub_o_hsize_ddr_bus_gpv),
        .htrans_ddr_bus_gpv_s0         (ddr_sub_o_htrans_ddr_bus_gpv),
        .hwdata_ddr_bus_gpv_s0         (ddr_sub_o_hwdata_ddr_bus_gpv),
        .hwrite_ddr_bus_gpv_s0         (ddr_sub_o_hwrite_ddr_bus_gpv),
        .hrdata_ddr_bus_gpv_s0         (ddr_sub_i_hrdata_ddr_bus_gpv),
        .hreadyout_ddr_bus_gpv_s0      (ddr_sub_i_hreadyout_ddr_bus_gpv),
        .hresp_ddr_bus_gpv_s0          (ddr_sub_i_hresp_ddr_bus_gpv),
        .hselx_ddr_bus_gpv_s0          (1'h1),
        .hready_ddr_bus_gpv_s0         (ddr_sub_i_hreadyout_ddr_bus_gpv),
        .i_ddr_busclk                  (ddr_crm_o_mclk_omc),
        .i_ddr_busresetn               (ddr_crm_o_mrstn_omc),
        .i_main2ddrclk                 (ddr_crm_o_clk_main2ddr),
        .i_main2ddrresetn              (ddr_crm_o_rstn_main2ddr),
        .i_periclk                     (ddr_crm_o_clk_peri2ddr),
        .i_periresetn                  (ddr_crm_o_rstn_peri2ddr),
        .mainclk                       (ddr_crm_o_mclk_omc),
        .mainclk_r                     (ddr_crm_o_mclk_omc),
        .mainresetn                    (ddr_crm_o_mrstn_omc),
        .mainresetn_r                  (ddr_crm_o_mrstn_omc)
    );

    ddr_sub
        #(.IB(11), .DB(128))
    u_ddr_sub (
        .i_clk_ddr_ref                 (ddr_crm_o_clk_ddr_ref),
        .i_rstn_ddr_ref                (ddr_crm_o_rstn_ddr_ref),
        .i_clk_peri2ddr                (ddr_crm_o_clk_peri2ddr),
        .i_rstn_peri2ddr               (ddr_crm_o_rstn_peri2ddr),
        .i_clk_peri2omc                (ddr_crm_o_sclk_omc),
        .i_rstn_peri2omc               (ddr_crm_o_srstn_omc),
        .i_clk_peri2phy                (ddr_crm_o_sclk_ddr_phy),
        .i_rstn_peri2phy               (ddr_crm_o_srstn_ddr_phy),
        .i_clk_ddr_phy                 (ddr_crm_o_mclk_ddr_phy),
        .i_rstn_ddr_phy                (ddr_crm_o_mrstn_ddr_phy),
        .i_clk_ddr_phym                (ddr_crm_o_clk_ddr_phym),
        .i_clk_ddr_omc                 (ddr_crm_o_mclk_omc),
        .i_rstn_ddr_omc                (ddr_crm_o_mrstn_omc),
        .o_clk_dfi                     (ddr_sub_o_clk_dfi),
        .i_psel_ddr_m0_deco            (i_psel_ddr_m0_deco),
        .i_penable_ddr_m0_deco         (i_penable_ddr_m0_deco),
        .i_paddr_ddr_m0_deco           (i_paddr_ddr_m0_deco),
        .i_pwrite_ddr_m0_deco          (i_pwrite_ddr_m0_deco),
        .i_pwdata_ddr_m0_deco          (i_pwdata_ddr_m0_deco),
        .o_prdata_ddr_m0_deco          (o_prdata_ddr_m0_deco),
        .o_pready_ddr_m0_deco          (o_pready_ddr_m0_deco),
        .o_pslverr_ddr_m0_deco         (o_pslverr_ddr_m0_deco),
        .o_psel_ddr_crm                (ddr_sub_o_psel_ddr_crm),
        .o_penable_ddr_crm             (ddr_sub_o_penable_ddr_crm),
        .o_paddr_ddr_crm               (ddr_sub_o_paddr_ddr_crm),
        .o_pwrite_ddr_crm              (ddr_sub_o_pwrite_ddr_crm),
        .o_pwdata_ddr_crm              (ddr_sub_o_pwdata_ddr_crm),
        .i_prdata_ddr_crm              (ddr_sub_i_prdata_ddr_crm),
        .o_haddr_ddr_bus_gpv           (ddr_sub_o_haddr_ddr_bus_gpv),
        .o_hburst_ddr_bus_gpv          (ddr_sub_o_hburst_ddr_bus_gpv),
        .o_hsize_ddr_bus_gpv           (ddr_sub_o_hsize_ddr_bus_gpv),
        .o_htrans_ddr_bus_gpv          (ddr_sub_o_htrans_ddr_bus_gpv),
        .o_hwdata_ddr_bus_gpv          (ddr_sub_o_hwdata_ddr_bus_gpv),
        .o_hwrite_ddr_bus_gpv          (ddr_sub_o_hwrite_ddr_bus_gpv),
        .i_hrdata_ddr_bus_gpv          (ddr_sub_i_hrdata_ddr_bus_gpv),
        .i_hreadyout_ddr_bus_gpv       (ddr_sub_i_hreadyout_ddr_bus_gpv),
        .i_hresp_ddr_bus_gpv           (ddr_sub_i_hresp_ddr_bus_gpv),
        .i_awid                        (ddr_bus_awid_ddr_m0),
        .i_awaddr                      (ddr_bus_awaddr_ddr_m0),
        .i_awlen                       (ddr_bus_awlen_ddr_m0),
        .i_awsize                      (ddr_bus_awsize_ddr_m0),
        .i_awburst                     (ddr_bus_awburst_ddr_m0),
        .i_awlock                      (ddr_bus_awlock_ddr_m0),
        .i_awcache                     (ddr_bus_awcache_ddr_m0),
        .i_awprot                      (ddr_bus_awprot_ddr_m0),
        .i_awvalid                     (ddr_bus_awvalid_ddr_m0),
        .o_awready                     (ddr_bus_awready_ddr_m0),
        .i_wdata                       (ddr_bus_wdata_ddr_m0),
        .i_wstrb                       (ddr_bus_wstrb_ddr_m0),
        .i_wlast                       (ddr_bus_wlast_ddr_m0),
        .i_wvalid                      (ddr_bus_wvalid_ddr_m0),
        .o_wready                      (ddr_bus_wready_ddr_m0),
        .o_bid                         (ddr_bus_bid_ddr_m0),
        .o_bresp                       (ddr_bus_bresp_ddr_m0),
        .o_bvalid                      (ddr_bus_bvalid_ddr_m0),
        .i_bready                      (ddr_bus_bready_ddr_m0),
        .i_arid                        (ddr_bus_arid_ddr_m0),
        .i_araddr                      (ddr_bus_araddr_ddr_m0),
        .i_arlen                       (ddr_bus_arlen_ddr_m0),
        .i_arsize                      (ddr_bus_arsize_ddr_m0),
        .i_arburst                     (ddr_bus_arburst_ddr_m0),
        .i_arlock                      (ddr_bus_arlock_ddr_m0),
        .i_arcache                     (ddr_bus_arcache_ddr_m0),
        .i_arprot                      (ddr_bus_arprot_ddr_m0),
        .i_arvalid                     (ddr_bus_arvalid_ddr_m0),
        .o_arready                     (ddr_bus_arready_ddr_m0),
        .o_rid                         (ddr_bus_rid_ddr_m0),
        .o_rdata                       (ddr_bus_rdata_ddr_m0),
        .o_rresp                       (ddr_bus_rresp_ddr_m0),
        .o_rlast                       (ddr_bus_rlast_ddr_m0),
        .o_rvalid                      (ddr_bus_rvalid_ddr_m0),
        .i_rready                      (ddr_bus_rready_ddr_m0),
        .o_irq_asp                     (o_irq_asp),
        .o_irq_overtemp                (o_irq_overtemp),
        .o_irq_hightemp                (o_irq_hightemp),
        .o_irq_cooldown                (o_irq_cooldown),
        .DDR_VREF0                     (DDR_VREF0),
        .DDR_VREF1                     (DDR_VREF1),
        .DDR_MEM_CKEIN                 (DDR_MEM_CKEIN),
        .DDR_MEM_CK_P                  (DDR_MEM_CK_P),
        .DDR_MEM_CK_N                  (DDR_MEM_CK_N),
        .DDR_MEM_CKE                   (DDR_MEM_CKE),
        .DDR_MEM_RESET_N               (DDR_MEM_RESET_N),
        .DDR_MEM_ODT                   (DDR_MEM_ODT),
        .DDR_MEM_CSN                   (DDR_MEM_CSN),
        .DDR_MEM_RASN                  (DDR_MEM_RASN),
        .DDR_MEM_CASN                  (DDR_MEM_CASN),
        .DDR_MEM_WEN                   (DDR_MEM_WEN),
        .DDR_MEM_BA                    (DDR_MEM_BA),
        .DDR_MEM_A                     (DDR_MEM_A),
        .DDR_MEM_DQ                    (DDR_MEM_DQ),
        .DDR_MEM_DM                    (DDR_MEM_DM),
        .DDR_MEM_DQS_P                 (DDR_MEM_DQS_P),
        .DDR_MEM_DQS_N                 (DDR_MEM_DQS_N),
        .DDR_ZQ                        (DDR_ZQ),
        .i_mode_phy_y                  (t_ddr_phy_phy_y),
        .i_mode_scan_y                 (t_ddr_phy_scan_y),
        .i_mode_nand_y                 (t_ddr_phy_nand_y),
        .i_mode_run_y                  (t_ddr_phy_run_y),
        .i_mode_mux_y                  (t_ddr_phy_mux_y),
        .i_mode_highz_y                (t_ddr_phy_highz_y),
        .i_test_ext_en_y               (t_ddr_phy_ext_en_y),
        .i_test_ext_out_y              (t_ddr_phy_ext_out_y),
        .i_test_ext_read_y             (t_ddr_phy_ext_read_y),
        .i_test_ext_cmosrcv_y          (t_ddr_phy_ext_cmosrcv_y),
        .i_test_ext_zq_force_y         (t_ddr_phy_ext_zq_force_y),
        .i_test_ext_zq_force_impp_y    (t_ddr_phy_ext_zq_force_impp_y),
        .i_test_ext_zq_force_impn_y    (t_ddr_phy_ext_zq_force_impn_y),
        .i_test_ext_zq_mode_dds_y      (t_ddr_phy_ext_zq_mode_dds_y),
        .i_test_ext_dfdqs_y            (t_ddr_phy_ext_dfdqs_y),
        .i_test_ext_ref_y              (t_ddr_phy_ext_ref_y),
        .i_test_ext_offsetc_y          (t_ddr_phy_ext_offsetc_y),
        .i_test_ext_rdlvl_en_y         (t_ddr_phy_ext_rdlvl_en_y),
        .i_test_ext_rdlvl_wr_en_y      (t_ddr_phy_ext_rdlvl_wr_en_y),
        .i_test_ext_gatelvl_en_y       (t_ddr_phy_ext_gatelvl_en_y),
        .i_test_ext_write_lvl_en_y     (t_ddr_phy_ext_write_lvl_en_y),
        .i_test_ext_ca_cal_en_y        (t_ddr_phy_ext_ca_cal_en_y),
        .i_test_ext_mode_y             (t_ddr_phy_ext_mode_y),
        .i_test_start_y                (t_ddr_phy_start_y),
        .i_test_ext_rdlvl_incr_adj_y   (t_ddr_phy_ext_rdlvl_incr_adj_y),
        .o_test_ctrl_div_out_400_a     (t_ddr_phy_ctrl_div_out_400_a),
        .o_test_ctrl_div_out_800_a     (t_ddr_phy_ctrl_div_out_800_a),
        .o_test_ext_zq_end_a           (t_ddr_phy_ext_zq_end_a),
        .o_test_ext_lock_value_a       (t_ddr_phy_ext_lock_value_a),
        .o_test_ext_clock_a            (t_ddr_phy_ext_clock_a),
        .o_test_ext_flock_a            (t_ddr_phy_ext_flock_a),
        .o_test_ext_locked_a           (t_ddr_phy_ext_locked_a),
        .o_test_ext_init_complete_a    (t_ddr_phy_ext_init_complete_a),
        .o_test_ext_rdlvl_vwmc_a       (t_ddr_phy_ext_rdlvl_vwmc_a),
        .o_test_err_a                  (t_ddr_phy_err_a),
        .o_test_oky_a                  (t_ddr_phy_oky_a),
        .test_se                       (test_se),
        .test_si                       (test_si),
        .test_so                       (test_so)
    );

endmodule