module main_crm (
    input           i_xtal         ,
    input           i_reset        ,
    output          o_cpu_aclk     ,
    output          o_cpu_areset   ,
    output          o_cpu_pclk     ,
    output          o_cpu_preset   ,
    output          o_peri_aclk    ,
    output          o_peri_areset  ,
    output          o_peri_pclk    ,
    output          o_peri_preset
);

endmodule