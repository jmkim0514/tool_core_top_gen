//==============================================================================
//
// Project : MVP
//
// Verilog RTL(Behavioral) model
//
// This confidential and proprietary source code may be used only as authorized
// by a licensing agreement from ALPHAHOLDINGS Limited. The entire notice above
// must be reproduced on all authorized copies and copies may only be made to
// the extent permitted by a licensing agreement from ALPHAHOLDINGS Limited.
//
// COPYRIGHT (C) ALPHAHOLDINGS, inc. 2022
//
//==============================================================================
// File name : mvp_hpdf
// Version : v1.1
// Description :
// Simulator : NC Verilog
// Created by : bhoh
// Date : 2023-08-28  15:48
//==============================================================================

module mvp_hpdf (
    input              i_rstn_cpu2mvp,
    input              i_clk_cpu2mvp,
    input              i_clk_xtal_y,
    input              i_clk_mvp2main,
    input              i_clk_dvp0_y,
    input              i_clk_dvp1_y,
    input              i_clk_dvp2_y,
    input              i_clk_dvp3_y,
    input              i_clk_dvp4_y,
    input              i_clk_dvp5_y,
    input              i_clk_dvp6_y,
    input              i_clk_dvp7_y,
    input              i_crm_test_mode,
    input              i_test_rstn,
    input              i_test_clk100,
    input              i_test_clk24,
    input              i_test_clk300,
    input              i_test_mode,
    input   [  5:  0]  t_tg_pll_p,
    input   [  9:  0]  t_tg_pll_m,
    input   [  2:  0]  t_tg_pll_s,
    input   [  1:  0]  t_tg_pll_lock_con_in,
    input   [  1:  0]  t_tg_pll_lock_con_out,
    input   [  1:  0]  t_tg_pll_lock_con_dly,
    input   [  1:  0]  t_tg_pll_lock_con_rev,
    input   [  4:  0]  t_tg_pll_tst_afc,
    input   [  1:  0]  t_tg_pll_icp,
    input              t_tg_pll_fin,
    input              t_tg_pll_resetb,
    input              t_tg_pll_bypass,
    input              t_tg_pll_tst_en,
    input              t_tg_pll_fsel,
    input              t_tg_pll_feed_en,
    input              t_tg_pll_lock_en,
    input              t_tg_pll_afcini_sel,
    input              t_tg_pll_vcoini_en,
    input              t_tg_pll_fout_mask,
    input              t_tg_pll_pbias_ctrl,
    input              t_tg_pll_pbias_ctrl_en,
    output             t_tg_pll_feed_out,
    output             t_tg_pll_lock,
    output             t_tg_pll_fout,
    output             t_tg_pll_sync_m_clk_out,
    output  [  4:  0]  t_tg_pll_afc_code,
    input   [  5:  0]  t_isp0_pll_p,
    input   [  9:  0]  t_isp0_pll_m,
    input   [  2:  0]  t_isp0_pll_s,
    input   [  1:  0]  t_isp0_pll_lock_con_in,
    input   [  1:  0]  t_isp0_pll_lock_con_out,
    input   [  1:  0]  t_isp0_pll_lock_con_dly,
    input   [  1:  0]  t_isp0_pll_lock_con_rev,
    input   [  4:  0]  t_isp0_pll_tst_afc,
    input   [  1:  0]  t_isp0_pll_icp,
    input              t_isp0_pll_fin,
    input              t_isp0_pll_resetb,
    input              t_isp0_pll_bypass,
    input              t_isp0_pll_tst_en,
    input              t_isp0_pll_fsel,
    input              t_isp0_pll_feed_en,
    input              t_isp0_pll_lock_en,
    input              t_isp0_pll_afcini_sel,
    input              t_isp0_pll_vcoini_en,
    input              t_isp0_pll_fout_mask,
    input              t_isp0_pll_pbias_ctrl,
    input              t_isp0_pll_pbias_ctrl_en,
    output             t_isp0_pll_feed_out,
    output             t_isp0_pll_lock,
    output             t_isp0_pll_fout,
    output             t_isp0_pll_sync_m_clk_out,
    output  [  4:  0]  t_isp0_pll_afc_code,
    input   [  5:  0]  t_isp1_pll_p,
    input   [  9:  0]  t_isp1_pll_m,
    input   [  2:  0]  t_isp1_pll_s,
    input   [  1:  0]  t_isp1_pll_lock_con_in,
    input   [  1:  0]  t_isp1_pll_lock_con_out,
    input   [  1:  0]  t_isp1_pll_lock_con_dly,
    input   [  1:  0]  t_isp1_pll_lock_con_rev,
    input   [  4:  0]  t_isp1_pll_tst_afc,
    input   [  1:  0]  t_isp1_pll_icp,
    input              t_isp1_pll_fin,
    input              t_isp1_pll_resetb,
    input              t_isp1_pll_bypass,
    input              t_isp1_pll_tst_en,
    input              t_isp1_pll_fsel,
    input              t_isp1_pll_feed_en,
    input              t_isp1_pll_lock_en,
    input              t_isp1_pll_afcini_sel,
    input              t_isp1_pll_vcoini_en,
    input              t_isp1_pll_fout_mask,
    input              t_isp1_pll_pbias_ctrl,
    input              t_isp1_pll_pbias_ctrl_en,
    output             t_isp1_pll_feed_out,
    output             t_isp1_pll_lock,
    output             t_isp1_pll_fout,
    output             t_isp1_pll_sync_m_clk_out,
    output  [  4:  0]  t_isp1_pll_afc_code,
    output             o_irq_wdma_err_00,
    output             o_irq_wdma_err_01,
    output             o_irq_wdma_err_02,
    output             o_irq_wdma_err_03,
    output             o_irq_wdma_err_04,
    output             o_irq_wdma_err_05,
    output             o_irq_wdma_err_06,
    output             o_irq_wdma_err_07,
    output             o_irq_wdma_done_00,
    output             o_irq_wdma_done_01,
    output             o_irq_wdma_done_02,
    output             o_irq_wdma_done_03,
    output             o_irq_wdma_done_04,
    output             o_irq_wdma_done_05,
    output             o_irq_wdma_done_06,
    output             o_irq_wdma_done_07,
    output             o_irq_rdma_err,
    output             o_irq_rdma_done,
    output             o_irq_rwdma_err,
    output             o_irq_gwdma_err,
    output             o_irq_bwdma_err,
    output             o_irq_rwdma_done,
    output             o_irq_gwdma_done,
    output             o_irq_bwdma_done,
    output             o_irq_qisp0_0,
    output             o_irq_qisp0_1,
    output             o_irq_qisp1_0,
    output             o_irq_qisp1_1,
    input              i_isp0_cis_dvp_v_y,
    input              i_isp0_cis_dvp_h_y,
    input              i_isp0_cis_dvp_pv_y,
    input   [  9:  0]  i_isp0_cis_dvp_p_y,
    input              i_isp1_cis_dvp_v_y,
    input              i_isp1_cis_dvp_h_y,
    input              i_isp1_cis_dvp_pv_y,
    input   [  9:  0]  i_isp1_cis_dvp_p_y,
    input              i_isp2_cis_dvp_v_y,
    input              i_isp2_cis_dvp_h_y,
    input              i_isp2_cis_dvp_pv_y,
    input   [  9:  0]  i_isp2_cis_dvp_p_y,
    input              i_isp3_cis_dvp_v_y,
    input              i_isp3_cis_dvp_h_y,
    input              i_isp3_cis_dvp_pv_y,
    input   [  9:  0]  i_isp3_cis_dvp_p_y,
    input              i_isp4_cis_dvp_v_y,
    input              i_isp4_cis_dvp_h_y,
    input              i_isp4_cis_dvp_pv_y,
    input   [  9:  0]  i_isp4_cis_dvp_p_y,
    input              i_isp5_cis_dvp_v_y,
    input              i_isp5_cis_dvp_h_y,
    input              i_isp5_cis_dvp_pv_y,
    input   [  9:  0]  i_isp5_cis_dvp_p_y,
    input              i_isp6_cis_dvp_v_y,
    input              i_isp6_cis_dvp_h_y,
    input              i_isp6_cis_dvp_pv_y,
    input   [  9:  0]  i_isp6_cis_dvp_p_y,
    input              i_isp7_cis_dvp_v_y,
    input              i_isp7_cis_dvp_h_y,
    input              i_isp7_cis_dvp_pv_y,
    input   [  9:  0]  i_isp7_cis_dvp_p_y,
    input   [ 38:  0]  i_ema,
    output             o_isp0_i2cm_scl_a,
    output             o_isp0_i2cm_sda_a,
    output             o_isp0_i2cm_sda_oe,
    input              i_isp0_i2cm_sda_y,
    output             o_isp1_i2cm_scl_a,
    output             o_isp1_i2cm_sda_a,
    output             o_isp1_i2cm_sda_oe,
    input              i_isp1_i2cm_sda_y,
    output             o_isp2_i2cm_scl_a,
    output             o_isp2_i2cm_sda_a,
    output             o_isp2_i2cm_sda_oe,
    input              i_isp2_i2cm_sda_y,
    output             o_isp3_i2cm_scl_a,
    output             o_isp3_i2cm_sda_a,
    output             o_isp3_i2cm_sda_oe,
    input              i_isp3_i2cm_sda_y,
    output             o_isp4_i2cm_scl_a,
    output             o_isp4_i2cm_sda_a,
    output             o_isp4_i2cm_sda_oe,
    input              i_isp4_i2cm_sda_y,
    output             o_isp5_i2cm_scl_a,
    output             o_isp5_i2cm_sda_a,
    output             o_isp5_i2cm_sda_oe,
    input              i_isp5_i2cm_sda_y,
    output             o_isp6_i2cm_scl_a,
    output             o_isp6_i2cm_sda_a,
    output             o_isp6_i2cm_sda_oe,
    input              i_isp6_i2cm_sda_y,
    output             o_isp7_i2cm_scl_a,
    output             o_isp7_i2cm_sda_a,
    output             o_isp7_i2cm_sda_oe,
    input              i_isp7_i2cm_sda_y,
    input              i_i2cs_scl_y,
    output             o_i2cs_sda_a,
    output             o_i2cs_sda_oe,
    input              i_i2cs_sda_y,
    output  [  9:  0]  o_isp0_cis_dvp_p_oe,
    output  [  9:  0]  o_isp1_cis_dvp_p_oe,
    output  [  9:  0]  o_isp2_cis_dvp_p_oe,
    output  [  9:  0]  o_isp3_cis_dvp_p_oe,
    output  [  9:  0]  o_isp4_cis_dvp_p_oe,
    output  [  9:  0]  o_isp5_cis_dvp_p_oe,
    output  [  9:  0]  o_isp6_cis_dvp_p_oe,
    output  [  9:  0]  o_isp7_cis_dvp_p_oe,
    output  [  9:  0]  o_isp0_cis_dvp_p_a,
    output  [  9:  0]  o_isp1_cis_dvp_p_a,
    output  [  9:  0]  o_isp2_cis_dvp_p_a,
    output  [  9:  0]  o_isp3_cis_dvp_p_a,
    output  [  9:  0]  o_isp4_cis_dvp_p_a,
    output  [  9:  0]  o_isp5_cis_dvp_p_a,
    output  [  9:  0]  o_isp6_cis_dvp_p_a,
    output  [  9:  0]  o_isp7_cis_dvp_p_a,
    output             o_tgclk_a,
    output             o_tg_dvp_v_a,
    output             o_tg_dvp_h_a,
    output  [ 31:  0]  o_tg_dvp_p_a,
    input              MIPI_CLKP_RX0,
    input              MIPI_CLKN_RX0,
    input   [  3:  0]  MIPI_DP_RX0,
    input   [  3:  0]  MIPI_DN_RX0,
    input              MIPI_CLKP_RX1,
    input              MIPI_CLKN_RX1,
    input   [  3:  0]  MIPI_DP_RX1,
    input   [  3:  0]  MIPI_DN_RX1,
    input              MIPI_CLKP_RX2,
    input              MIPI_CLKN_RX2,
    input   [  3:  0]  MIPI_DP_RX2,
    input   [  3:  0]  MIPI_DN_RX2,
    input              MIPI_CLKP_RX3,
    input              MIPI_CLKN_RX3,
    input   [  3:  0]  MIPI_DP_RX3,
    input   [  3:  0]  MIPI_DN_RX3,
    input              MIPI_CHIP_EN_MR0,
    output             MIPI_HS_CKO_RX0,
    output  [  3:  0]  MIPI_HS_DO_RX0,
    output             MIPI_TEST_VMON_OUT_RX0,
    input              MIPI_CLKP_RX4,
    input              MIPI_CLKN_RX4,
    input   [  3:  0]  MIPI_DP_RX4,
    input   [  3:  0]  MIPI_DN_RX4,
    input              MIPI_CLKP_RX5,
    input              MIPI_CLKN_RX5,
    input   [  3:  0]  MIPI_DP_RX5,
    input   [  3:  0]  MIPI_DN_RX5,
    input              MIPI_CLKP_RX6,
    input              MIPI_CLKN_RX6,
    input   [  3:  0]  MIPI_DP_RX6,
    input   [  3:  0]  MIPI_DN_RX6,
    input              MIPI_CLKP_RX7,
    input              MIPI_CLKN_RX7,
    input   [  3:  0]  MIPI_DP_RX7,
    input   [  3:  0]  MIPI_DN_RX7,
    input              MIPI_CHIP_EN_MR1,
    output             MIPI_HS_CKO_RX4,
    output  [  3:  0]  MIPI_HS_DO_RX4,
    output             MIPI_TEST_VMON_OUT_RX4,
    input              MIPI_CHIP_EN_TX,
    output             MIPI_CLKP_TX,
    output             MIPI_CLKN_TX,
    output  [  3:  0]  MIPI_DP_TX,
    output  [  3:  0]  MIPI_DN_TX,
    output             MIPI_HS_CKO_TX,
    output  [  3:  0]  MIPI_HS_DO_TX,
    output             MIPI_TEST_VMON_OUT_TX,
    output             MIPI_TEST_CLK_A0,
    input              i_psel_cpu2mvp,
    input              i_penable_cpu2mvp,
    input              i_pwrite_cpu2mvp,
    input   [ 31:  0]  i_paddr_cpu2mvp,
    input   [ 31:  0]  i_pwdata_cpu2mvp,
    output             o_pready_cpu2mvp,
    output  [ 31:  0]  o_prdata_cpu2mvp,
    output             o_pslverr_cpu2mvp,
    output  [  1:  0]  o_awid_rgb2main,
    output             o_awvalid_rgb2main,
    input              i_awready_rgb2main,
    output  [ 31:  0]  o_awaddr_rgb2main,
    output  [  2:  0]  o_awprot_rgb2main,
    output  [  7:  0]  o_awlen_rgb2main,
    output  [  2:  0]  o_awsize_rgb2main,
    output  [  1:  0]  o_awburst_rgb2main,
    output             o_awlock_rgb2main,
    output  [  3:  0]  o_awcache_rgb2main,
    output             o_wvalid_rgb2main,
    input              i_wready_rgb2main,
    output  [127:  0]  o_wdata_rgb2main,
    output  [ 15:  0]  o_wstrb_rgb2main,
    output             o_wlast_rgb2main,
    input   [  1:  0]  i_bid_rgb2main,
    input              i_bvalid_rgb2main,
    output             o_bready_rgb2main,
    input   [  1:  0]  i_bresp_rgb2main,
    output  [  1:  0]  o_arid_rgb2main,
    output  [  2:  0]  o_arprot_rgb2main,
    output             o_arvalid_rgb2main,
    input              i_arready_rgb2main,
    output  [ 31:  0]  o_araddr_rgb2main,
    output  [  7:  0]  o_arlen_rgb2main,
    output  [  2:  0]  o_arsize_rgb2main,
    output  [  1:  0]  o_arburst_rgb2main,
    output             o_arlock_rgb2main,
    output  [  3:  0]  o_arcache_rgb2main,
    input              i_rvalid_rgb2main,
    input   [  1:  0]  i_rid_rgb2main,
    output             o_rready_rgb2main,
    input   [127:  0]  i_rdata_rgb2main,
    input              i_rlast_rgb2main,
    input   [  1:  0]  i_rresp_rgb2main,
    output  [  1:  0]  o_awuser_rgb2main,
    output  [  1:  0]  o_aruser_rgb2main,
    output  [  1:  0]  o_awid_isp2main_0,
    output             o_awvalid_isp2main_0,
    input              i_awready_isp2main_0,
    output  [ 31:  0]  o_awaddr_isp2main_0,
    output  [  2:  0]  o_awprot_isp2main_0,
    output  [  7:  0]  o_awlen_isp2main_0,
    output  [  2:  0]  o_awsize_isp2main_0,
    output  [  1:  0]  o_awburst_isp2main_0,
    output             o_awlock_isp2main_0,
    output  [  3:  0]  o_awcache_isp2main_0,
    output             o_wvalid_isp2main_0,
    input              i_wready_isp2main_0,
    output  [127:  0]  o_wdata_isp2main_0,
    output  [ 15:  0]  o_wstrb_isp2main_0,
    output             o_wlast_isp2main_0,
    input   [  1:  0]  i_bid_isp2main_0,
    input              i_bvalid_isp2main_0,
    output             o_bready_isp2main_0,
    input   [  1:  0]  i_bresp_isp2main_0,
    output  [  1:  0]  o_arid_isp2main_0,
    output  [  2:  0]  o_arprot_isp2main_0,
    output             o_arvalid_isp2main_0,
    input              i_arready_isp2main_0,
    output  [ 31:  0]  o_araddr_isp2main_0,
    output  [  7:  0]  o_arlen_isp2main_0,
    output  [  2:  0]  o_arsize_isp2main_0,
    output  [  1:  0]  o_arburst_isp2main_0,
    output             o_arlock_isp2main_0,
    output  [  3:  0]  o_arcache_isp2main_0,
    input   [  1:  0]  i_rid_isp2main_0,
    input              i_rvalid_isp2main_0,
    output             o_rready_isp2main_0,
    input   [127:  0]  i_rdata_isp2main_0,
    input              i_rlast_isp2main_0,
    input   [  1:  0]  i_rresp_isp2main_0,
    output  [  1:  0]  o_awuser_isp2main_0,
    output  [  1:  0]  o_aruser_isp2main_0,
    output  [  1:  0]  o_awid_isp2main_1,
    output             o_awvalid_isp2main_1,
    input              i_awready_isp2main_1,
    output  [ 31:  0]  o_awaddr_isp2main_1,
    output  [  2:  0]  o_awprot_isp2main_1,
    output  [  7:  0]  o_awlen_isp2main_1,
    output  [  2:  0]  o_awsize_isp2main_1,
    output  [  1:  0]  o_awburst_isp2main_1,
    output             o_awlock_isp2main_1,
    output  [  3:  0]  o_awcache_isp2main_1,
    output             o_wvalid_isp2main_1,
    input              i_wready_isp2main_1,
    output  [127:  0]  o_wdata_isp2main_1,
    output  [ 15:  0]  o_wstrb_isp2main_1,
    output             o_wlast_isp2main_1,
    input   [  1:  0]  i_bid_isp2main_1,
    input              i_bvalid_isp2main_1,
    output             o_bready_isp2main_1,
    input   [  1:  0]  i_bresp_isp2main_1,
    output  [  1:  0]  o_arid_isp2main_1,
    output  [  2:  0]  o_arprot_isp2main_1,
    output             o_arvalid_isp2main_1,
    input              i_arready_isp2main_1,
    output  [ 31:  0]  o_araddr_isp2main_1,
    output  [  7:  0]  o_arlen_isp2main_1,
    output  [  2:  0]  o_arsize_isp2main_1,
    output  [  1:  0]  o_arburst_isp2main_1,
    output             o_arlock_isp2main_1,
    output  [  3:  0]  o_arcache_isp2main_1,
    input   [  1:  0]  i_rid_isp2main_1,
    input              i_rvalid_isp2main_1,
    output             o_rready_isp2main_1,
    input   [127:  0]  i_rdata_isp2main_1,
    input              i_rlast_isp2main_1,
    input   [  1:  0]  i_rresp_isp2main_1,
    output  [  1:  0]  o_awuser_isp2main_1,
    output  [  1:  0]  o_aruser_isp2main_1
);

    wire            mvp_crm_o_pll_tg_norm_resetb;
    wire            mvp_crm_o_pll_tg_norm_bypass;
    wire    [ 5:0]  mvp_crm_o_pll_tg_norm_p;
    wire    [ 9:0]  mvp_crm_o_pll_tg_norm_m;
    wire    [ 2:0]  mvp_crm_o_pll_tg_norm_s;
    wire            mvp_crm_o_pll_tg_norm_lock_en;
    wire    [ 1:0]  mvp_crm_o_pll_tg_norm_lock_con_in;
    wire    [ 1:0]  mvp_crm_o_pll_tg_norm_lock_con_out;
    wire    [ 1:0]  mvp_crm_o_pll_tg_norm_lock_con_dly;
    wire    [ 1:0]  mvp_crm_o_pll_tg_norm_lock_con_rev;
    wire            mvp_crm_o_pll_tg_norm_feed_en;
    wire            mvp_crm_o_pll_tg_norm_fsel;
    wire            mvp_crm_o_pll_tg_norm_tst_en;
    wire    [ 4:0]  mvp_crm_o_pll_tg_norm_tst_afc;
    wire            mvp_crm_o_pll_tg_norm_afcini_sel;
    wire            mvp_crm_o_pll_tg_norm_vcoini_en;
    wire            mvp_crm_o_pll_tg_norm_fout_mask;
    wire            mvp_crm_o_pll_tg_norm_pbias_ctrl;
    wire            mvp_crm_o_pll_tg_norm_pbias_ctrl_en;
    wire    [ 1:0]  mvp_crm_o_pll_tg_norm_icp;
    wire            mvp_crm_o_pll_isp0_norm_resetb;
    wire            mvp_crm_o_pll_isp0_norm_bypass;
    wire    [ 5:0]  mvp_crm_o_pll_isp0_norm_p;
    wire    [ 9:0]  mvp_crm_o_pll_isp0_norm_m;
    wire    [ 2:0]  mvp_crm_o_pll_isp0_norm_s;
    wire            mvp_crm_o_pll_isp0_norm_lock_en;
    wire    [ 1:0]  mvp_crm_o_pll_isp0_norm_lock_con_in;
    wire    [ 1:0]  mvp_crm_o_pll_isp0_norm_lock_con_out;
    wire    [ 1:0]  mvp_crm_o_pll_isp0_norm_lock_con_dly;
    wire    [ 1:0]  mvp_crm_o_pll_isp0_norm_lock_con_rev;
    wire            mvp_crm_o_pll_isp0_norm_feed_en;
    wire            mvp_crm_o_pll_isp0_norm_fsel;
    wire            mvp_crm_o_pll_isp0_norm_tst_en;
    wire    [ 4:0]  mvp_crm_o_pll_isp0_norm_tst_afc;
    wire            mvp_crm_o_pll_isp0_norm_afcini_sel;
    wire            mvp_crm_o_pll_isp0_norm_vcoini_en;
    wire            mvp_crm_o_pll_isp0_norm_fout_mask;
    wire            mvp_crm_o_pll_isp0_norm_pbias_ctrl;
    wire            mvp_crm_o_pll_isp0_norm_pbias_ctrl_en;
    wire    [ 1:0]  mvp_crm_o_pll_isp0_norm_icp;
    wire            mvp_crm_o_pll_isp1_norm_resetb;
    wire            mvp_crm_o_pll_isp1_norm_bypass;
    wire    [ 5:0]  mvp_crm_o_pll_isp1_norm_p;
    wire    [ 9:0]  mvp_crm_o_pll_isp1_norm_m;
    wire    [ 2:0]  mvp_crm_o_pll_isp1_norm_s;
    wire            mvp_crm_o_pll_isp1_norm_lock_en;
    wire    [ 1:0]  mvp_crm_o_pll_isp1_norm_lock_con_in;
    wire    [ 1:0]  mvp_crm_o_pll_isp1_norm_lock_con_out;
    wire    [ 1:0]  mvp_crm_o_pll_isp1_norm_lock_con_dly;
    wire    [ 1:0]  mvp_crm_o_pll_isp1_norm_lock_con_rev;
    wire            mvp_crm_o_pll_isp1_norm_feed_en;
    wire            mvp_crm_o_pll_isp1_norm_fsel;
    wire            mvp_crm_o_pll_isp1_norm_tst_en;
    wire    [ 4:0]  mvp_crm_o_pll_isp1_norm_tst_afc;
    wire            mvp_crm_o_pll_isp1_norm_afcini_sel;
    wire            mvp_crm_o_pll_isp1_norm_vcoini_en;
    wire            mvp_crm_o_pll_isp1_norm_fout_mask;
    wire            mvp_crm_o_pll_isp1_norm_pbias_ctrl;
    wire            mvp_crm_o_pll_isp1_norm_pbias_ctrl_en;
    wire    [ 1:0]  mvp_crm_o_pll_isp1_norm_icp;
    wire            mvp_crm_o_clk_phy_ref;
    wire            mvp_crm_o_clk_riscv_timer0;
    wire            mvp_crm_o_rstn_riscv_timer0;
    wire            mvp_crm_o_clk_riscv_timer1;
    wire            mvp_crm_o_rstn_riscv_timer1;
    wire            mvp_crm_o_clk_cpu2mvp;
    wire            mvp_crm_o_rstn_cpu2mvp;
    wire            mvp_crm_o_sclk_wdma0;
    wire            mvp_crm_o_srstn_wdma0;
    wire            mvp_crm_o_sclk_wdma1;
    wire            mvp_crm_o_srstn_wdma1;
    wire            mvp_crm_o_sclk_wdma2;
    wire            mvp_crm_o_srstn_wdma2;
    wire            mvp_crm_o_sclk_wdma3;
    wire            mvp_crm_o_srstn_wdma3;
    wire            mvp_crm_o_sclk_wdma4;
    wire            mvp_crm_o_srstn_wdma4;
    wire            mvp_crm_o_sclk_wdma5;
    wire            mvp_crm_o_srstn_wdma5;
    wire            mvp_crm_o_sclk_wdma6;
    wire            mvp_crm_o_srstn_wdma6;
    wire            mvp_crm_o_sclk_wdma7;
    wire            mvp_crm_o_srstn_wdma7;
    wire            mvp_crm_o_sclk_y2r_dma;
    wire            mvp_crm_o_srstn_y2r_dma;
    wire            mvp_crm_o_sclk_rdma;
    wire            mvp_crm_o_srstn_rdma;
    wire            mvp_crm_o_clk_mvp2main;
    wire            mvp_crm_o_rstn_mvp2main;
    wire            mvp_crm_o_mclk_wdma0;
    wire            mvp_crm_o_mrstn_wdma0;
    wire            mvp_crm_o_mclk_wdma1;
    wire            mvp_crm_o_mrstn_wdma1;
    wire            mvp_crm_o_mclk_wdma2;
    wire            mvp_crm_o_mrstn_wdma2;
    wire            mvp_crm_o_mclk_wdma3;
    wire            mvp_crm_o_mrstn_wdma3;
    wire            mvp_crm_o_mclk_wdma4;
    wire            mvp_crm_o_mrstn_wdma4;
    wire            mvp_crm_o_mclk_wdma5;
    wire            mvp_crm_o_mrstn_wdma5;
    wire            mvp_crm_o_mclk_wdma6;
    wire            mvp_crm_o_mrstn_wdma6;
    wire            mvp_crm_o_mclk_wdma7;
    wire            mvp_crm_o_mrstn_wdma7;
    wire            mvp_crm_o_mclk_y2r_dma;
    wire            mvp_crm_o_mrstn_y2r_dma;
    wire            mvp_crm_o_clk_riscv;
    wire            mvp_crm_o_rstn_riscv;
    wire            mvp_crm_o_mclk_rdma;
    wire            mvp_crm_o_mrstn_rdma;
    wire            mvp_crm_o_clk_tg;
    wire            mvp_crm_o_rstn_tg;
    wire            mvp_crm_o_clk_yuv2rgb;
    wire            mvp_crm_o_rstn_yuv2rgb;
    wire            mvp_crm_o_clk_dvp0;
    wire            mvp_crm_o_rstn_dvp0;
    wire            mvp_crm_o_clk_dvp1;
    wire            mvp_crm_o_rstn_dvp1;
    wire            mvp_crm_o_clk_dvp2;
    wire            mvp_crm_o_rstn_dvp2;
    wire            mvp_crm_o_clk_dvp3;
    wire            mvp_crm_o_rstn_dvp3;
    wire            mvp_crm_o_clk_dvp4;
    wire            mvp_crm_o_rstn_dvp4;
    wire            mvp_crm_o_clk_dvp5;
    wire            mvp_crm_o_rstn_dvp5;
    wire            mvp_crm_o_clk_dvp6;
    wire            mvp_crm_o_rstn_dvp6;
    wire            mvp_crm_o_clk_dvp7;
    wire            mvp_crm_o_rstn_dvp7;
    wire            mvp_crm_o_clk_isp0_clk;
    wire            mvp_crm_o_rstn_isp0_clk;
    wire            mvp_crm_o_clk_isp1_clk;
    wire            mvp_crm_o_rstn_isp1_clk;
    wire            mvp_crm_o_clk_isp2_clk;
    wire            mvp_crm_o_rstn_isp2_clk;
    wire            mvp_crm_o_clk_isp3_clk;
    wire            mvp_crm_o_rstn_isp3_clk;
    wire            mvp_crm_o_clk_isp4_clk;
    wire            mvp_crm_o_rstn_isp4_clk;
    wire            mvp_crm_o_clk_isp5_clk;
    wire            mvp_crm_o_rstn_isp5_clk;
    wire            mvp_crm_o_clk_isp6_clk;
    wire            mvp_crm_o_rstn_isp6_clk;
    wire            mvp_crm_o_clk_isp7_clk;
    wire            mvp_crm_o_rstn_isp7_clk;
    wire            tg_pll_o_feed_out;
    wire            tg_pll_o_lock;
    wire            tg_pll_o_fout;
    wire            tg_pll_o_sync_m_clk_out;
    wire    [ 4:0]  tg_pll_o_afc_code;
    wire            isp0_pll_o_feed_out;
    wire            isp0_pll_o_lock;
    wire            isp0_pll_o_fout;
    wire            isp0_pll_o_sync_m_clk_out;
    wire    [ 4:0]  isp0_pll_o_afc_code;
    wire            isp1_pll_o_feed_out;
    wire            isp1_pll_o_lock;
    wire            isp1_pll_o_fout;
    wire            isp1_pll_o_sync_m_clk_out;
    wire    [ 4:0]  isp1_pll_o_afc_code;
    wire            mvp_sub_o_mvp_crm_psel;
    wire            mvp_sub_o_mvp_crm_penable;
    wire            mvp_sub_o_mvp_crm_pwrite;
    wire    [11:0]  mvp_sub_o_mvp_crm_paddr;
    wire    [31:0]  mvp_sub_o_mvp_crm_pwdata;
    wire    [31:0]  mvp_sub_i_mvp_crm_prdata;

    assign  t_isp0_pll_afc_code[4:0] = isp0_pll_o_afc_code[4:0];
    assign  t_isp0_pll_feed_out = isp0_pll_o_feed_out;
    assign  t_isp0_pll_fout = isp0_pll_o_fout;
    assign  t_isp0_pll_lock = isp0_pll_o_lock;
    assign  t_isp0_pll_sync_m_clk_out = isp0_pll_o_sync_m_clk_out;
    assign  t_isp1_pll_afc_code[4:0] = isp1_pll_o_afc_code[4:0];
    assign  t_isp1_pll_feed_out = isp1_pll_o_feed_out;
    assign  t_isp1_pll_fout = isp1_pll_o_fout;
    assign  t_isp1_pll_lock = isp1_pll_o_lock;
    assign  t_isp1_pll_sync_m_clk_out = isp1_pll_o_sync_m_clk_out;
    assign  t_tg_pll_afc_code[4:0] = tg_pll_o_afc_code[4:0];
    assign  t_tg_pll_feed_out = tg_pll_o_feed_out;
    assign  t_tg_pll_fout = tg_pll_o_fout;
    assign  t_tg_pll_lock = tg_pll_o_lock;
    assign  t_tg_pll_sync_m_clk_out = tg_pll_o_sync_m_clk_out;

    mvp_crm_mvp u_mvp_crm (
        .i_rstn_mvp                      (i_rstn_cpu2mvp),
        .i_apb_pclk                      (i_clk_cpu2mvp),
        .i_apb_prstn                     (i_rstn_cpu2mvp),
        .i_apb_psel                      (mvp_sub_o_mvp_crm_psel),
        .i_apb_penable                   (mvp_sub_o_mvp_crm_penable),
        .i_apb_pwrite                    (mvp_sub_o_mvp_crm_pwrite),
        .i_apb_paddr                     (mvp_sub_o_mvp_crm_paddr),
        .i_apb_pwdata                    (mvp_sub_o_mvp_crm_pwdata),
        .o_apb_prdata                    (mvp_sub_i_mvp_crm_prdata),
        .o_pll_tg_norm_resetb            (mvp_crm_o_pll_tg_norm_resetb),
        .o_pll_tg_norm_bypass            (mvp_crm_o_pll_tg_norm_bypass),
        .o_pll_tg_norm_p                 (mvp_crm_o_pll_tg_norm_p),
        .o_pll_tg_norm_m                 (mvp_crm_o_pll_tg_norm_m),
        .o_pll_tg_norm_s                 (mvp_crm_o_pll_tg_norm_s),
        .i_pll_tg_lock                   (tg_pll_o_lock),
        .i_pll_tg_feed_out               (tg_pll_o_feed_out),
        .i_pll_tg_sync_m_clk_out         (tg_pll_o_sync_m_clk_out),
        .i_pll_tg_afc_code               (tg_pll_o_afc_code),
        .o_pll_tg_norm_lock_en           (mvp_crm_o_pll_tg_norm_lock_en),
        .o_pll_tg_norm_lock_con_in       (mvp_crm_o_pll_tg_norm_lock_con_in),
        .o_pll_tg_norm_lock_con_out      (mvp_crm_o_pll_tg_norm_lock_con_out),
        .o_pll_tg_norm_lock_con_dly      (mvp_crm_o_pll_tg_norm_lock_con_dly),
        .o_pll_tg_norm_lock_con_rev      (mvp_crm_o_pll_tg_norm_lock_con_rev),
        .o_pll_tg_norm_feed_en           (mvp_crm_o_pll_tg_norm_feed_en),
        .o_pll_tg_norm_fsel              (mvp_crm_o_pll_tg_norm_fsel),
        .o_pll_tg_norm_tst_en            (mvp_crm_o_pll_tg_norm_tst_en),
        .o_pll_tg_norm_tst_afc           (mvp_crm_o_pll_tg_norm_tst_afc),
        .o_pll_tg_norm_afcini_sel        (mvp_crm_o_pll_tg_norm_afcini_sel),
        .o_pll_tg_norm_vcoini_en         (mvp_crm_o_pll_tg_norm_vcoini_en),
        .o_pll_tg_norm_fout_mask         (mvp_crm_o_pll_tg_norm_fout_mask),
        .o_pll_tg_norm_pbias_ctrl        (mvp_crm_o_pll_tg_norm_pbias_ctrl),
        .o_pll_tg_norm_pbias_ctrl_en     (mvp_crm_o_pll_tg_norm_pbias_ctrl_en),
        .o_pll_tg_norm_icp               (mvp_crm_o_pll_tg_norm_icp),
        .o_pll_isp0_norm_resetb          (mvp_crm_o_pll_isp0_norm_resetb),
        .o_pll_isp0_norm_bypass          (mvp_crm_o_pll_isp0_norm_bypass),
        .o_pll_isp0_norm_p               (mvp_crm_o_pll_isp0_norm_p),
        .o_pll_isp0_norm_m               (mvp_crm_o_pll_isp0_norm_m),
        .o_pll_isp0_norm_s               (mvp_crm_o_pll_isp0_norm_s),
        .i_pll_isp0_lock                 (isp0_pll_o_lock),
        .i_pll_isp0_feed_out             (isp0_pll_o_feed_out),
        .i_pll_isp0_sync_m_clk_out       (isp0_pll_o_sync_m_clk_out),
        .i_pll_isp0_afc_code             (isp0_pll_o_afc_code),
        .o_pll_isp0_norm_lock_en         (mvp_crm_o_pll_isp0_norm_lock_en),
        .o_pll_isp0_norm_lock_con_in     (mvp_crm_o_pll_isp0_norm_lock_con_in),
        .o_pll_isp0_norm_lock_con_out    (mvp_crm_o_pll_isp0_norm_lock_con_out),
        .o_pll_isp0_norm_lock_con_dly    (mvp_crm_o_pll_isp0_norm_lock_con_dly),
        .o_pll_isp0_norm_lock_con_rev    (mvp_crm_o_pll_isp0_norm_lock_con_rev),
        .o_pll_isp0_norm_feed_en         (mvp_crm_o_pll_isp0_norm_feed_en),
        .o_pll_isp0_norm_fsel            (mvp_crm_o_pll_isp0_norm_fsel),
        .o_pll_isp0_norm_tst_en          (mvp_crm_o_pll_isp0_norm_tst_en),
        .o_pll_isp0_norm_tst_afc         (mvp_crm_o_pll_isp0_norm_tst_afc),
        .o_pll_isp0_norm_afcini_sel      (mvp_crm_o_pll_isp0_norm_afcini_sel),
        .o_pll_isp0_norm_vcoini_en       (mvp_crm_o_pll_isp0_norm_vcoini_en),
        .o_pll_isp0_norm_fout_mask       (mvp_crm_o_pll_isp0_norm_fout_mask),
        .o_pll_isp0_norm_pbias_ctrl      (mvp_crm_o_pll_isp0_norm_pbias_ctrl),
        .o_pll_isp0_norm_pbias_ctrl_en   (mvp_crm_o_pll_isp0_norm_pbias_ctrl_en),
        .o_pll_isp0_norm_icp             (mvp_crm_o_pll_isp0_norm_icp),
        .o_pll_isp1_norm_resetb          (mvp_crm_o_pll_isp1_norm_resetb),
        .o_pll_isp1_norm_bypass          (mvp_crm_o_pll_isp1_norm_bypass),
        .o_pll_isp1_norm_p               (mvp_crm_o_pll_isp1_norm_p),
        .o_pll_isp1_norm_m               (mvp_crm_o_pll_isp1_norm_m),
        .o_pll_isp1_norm_s               (mvp_crm_o_pll_isp1_norm_s),
        .i_pll_isp1_lock                 (isp1_pll_o_lock),
        .i_pll_isp1_feed_out             (isp1_pll_o_feed_out),
        .i_pll_isp1_sync_m_clk_out       (isp1_pll_o_sync_m_clk_out),
        .i_pll_isp1_afc_code             (isp1_pll_o_afc_code),
        .o_pll_isp1_norm_lock_en         (mvp_crm_o_pll_isp1_norm_lock_en),
        .o_pll_isp1_norm_lock_con_in     (mvp_crm_o_pll_isp1_norm_lock_con_in),
        .o_pll_isp1_norm_lock_con_out    (mvp_crm_o_pll_isp1_norm_lock_con_out),
        .o_pll_isp1_norm_lock_con_dly    (mvp_crm_o_pll_isp1_norm_lock_con_dly),
        .o_pll_isp1_norm_lock_con_rev    (mvp_crm_o_pll_isp1_norm_lock_con_rev),
        .o_pll_isp1_norm_feed_en         (mvp_crm_o_pll_isp1_norm_feed_en),
        .o_pll_isp1_norm_fsel            (mvp_crm_o_pll_isp1_norm_fsel),
        .o_pll_isp1_norm_tst_en          (mvp_crm_o_pll_isp1_norm_tst_en),
        .o_pll_isp1_norm_tst_afc         (mvp_crm_o_pll_isp1_norm_tst_afc),
        .o_pll_isp1_norm_afcini_sel      (mvp_crm_o_pll_isp1_norm_afcini_sel),
        .o_pll_isp1_norm_vcoini_en       (mvp_crm_o_pll_isp1_norm_vcoini_en),
        .o_pll_isp1_norm_fout_mask       (mvp_crm_o_pll_isp1_norm_fout_mask),
        .o_pll_isp1_norm_pbias_ctrl      (mvp_crm_o_pll_isp1_norm_pbias_ctrl),
        .o_pll_isp1_norm_pbias_ctrl_en   (mvp_crm_o_pll_isp1_norm_pbias_ctrl_en),
        .o_pll_isp1_norm_icp             (mvp_crm_o_pll_isp1_norm_icp),
        .i_clk_xtal_y                    (i_clk_xtal_y),
        .i_clk_cpu2mvp                   (i_clk_cpu2mvp),
        .i_clk_mvp2main                  (i_clk_mvp2main),
        .i_pll_tg                        (tg_pll_o_fout),
        .i_clk_dvp0_y                    (i_clk_dvp0_y),
        .i_clk_dvp1_y                    (i_clk_dvp1_y),
        .i_clk_dvp2_y                    (i_clk_dvp2_y),
        .i_clk_dvp3_y                    (i_clk_dvp3_y),
        .i_clk_dvp4_y                    (i_clk_dvp4_y),
        .i_clk_dvp5_y                    (i_clk_dvp5_y),
        .i_clk_dvp6_y                    (i_clk_dvp6_y),
        .i_clk_dvp7_y                    (i_clk_dvp7_y),
        .i_pll_isp0                      (isp0_pll_o_fout),
        .i_pll_isp1                      (isp1_pll_o_fout),
        .o_clk_phy_ref                   (mvp_crm_o_clk_phy_ref),
        .o_clk_riscv_timer0              (mvp_crm_o_clk_riscv_timer0),
        .o_rstn_riscv_timer0             (mvp_crm_o_rstn_riscv_timer0),
        .o_clk_riscv_timer1              (mvp_crm_o_clk_riscv_timer1),
        .o_rstn_riscv_timer1             (mvp_crm_o_rstn_riscv_timer1),
        .o_clk_cpu2mvp                   (mvp_crm_o_clk_cpu2mvp),
        .o_rstn_cpu2mvp                  (mvp_crm_o_rstn_cpu2mvp),
        .o_sclk_wdma0                    (mvp_crm_o_sclk_wdma0),
        .o_srstn_wdma0                   (mvp_crm_o_srstn_wdma0),
        .o_sclk_wdma1                    (mvp_crm_o_sclk_wdma1),
        .o_srstn_wdma1                   (mvp_crm_o_srstn_wdma1),
        .o_sclk_wdma2                    (mvp_crm_o_sclk_wdma2),
        .o_srstn_wdma2                   (mvp_crm_o_srstn_wdma2),
        .o_sclk_wdma3                    (mvp_crm_o_sclk_wdma3),
        .o_srstn_wdma3                   (mvp_crm_o_srstn_wdma3),
        .o_sclk_wdma4                    (mvp_crm_o_sclk_wdma4),
        .o_srstn_wdma4                   (mvp_crm_o_srstn_wdma4),
        .o_sclk_wdma5                    (mvp_crm_o_sclk_wdma5),
        .o_srstn_wdma5                   (mvp_crm_o_srstn_wdma5),
        .o_sclk_wdma6                    (mvp_crm_o_sclk_wdma6),
        .o_srstn_wdma6                   (mvp_crm_o_srstn_wdma6),
        .o_sclk_wdma7                    (mvp_crm_o_sclk_wdma7),
        .o_srstn_wdma7                   (mvp_crm_o_srstn_wdma7),
        .o_sclk_y2r_dma                  (mvp_crm_o_sclk_y2r_dma),
        .o_srstn_y2r_dma                 (mvp_crm_o_srstn_y2r_dma),
        .o_sclk_rdma                     (mvp_crm_o_sclk_rdma),
        .o_srstn_rdma                    (mvp_crm_o_srstn_rdma),
        .o_clk_mvp2main                  (mvp_crm_o_clk_mvp2main),
        .o_rstn_mvp2main                 (mvp_crm_o_rstn_mvp2main),
        .o_mclk_wdma0                    (mvp_crm_o_mclk_wdma0),
        .o_mrstn_wdma0                   (mvp_crm_o_mrstn_wdma0),
        .o_mclk_wdma1                    (mvp_crm_o_mclk_wdma1),
        .o_mrstn_wdma1                   (mvp_crm_o_mrstn_wdma1),
        .o_mclk_wdma2                    (mvp_crm_o_mclk_wdma2),
        .o_mrstn_wdma2                   (mvp_crm_o_mrstn_wdma2),
        .o_mclk_wdma3                    (mvp_crm_o_mclk_wdma3),
        .o_mrstn_wdma3                   (mvp_crm_o_mrstn_wdma3),
        .o_mclk_wdma4                    (mvp_crm_o_mclk_wdma4),
        .o_mrstn_wdma4                   (mvp_crm_o_mrstn_wdma4),
        .o_mclk_wdma5                    (mvp_crm_o_mclk_wdma5),
        .o_mrstn_wdma5                   (mvp_crm_o_mrstn_wdma5),
        .o_mclk_wdma6                    (mvp_crm_o_mclk_wdma6),
        .o_mrstn_wdma6                   (mvp_crm_o_mrstn_wdma6),
        .o_mclk_wdma7                    (mvp_crm_o_mclk_wdma7),
        .o_mrstn_wdma7                   (mvp_crm_o_mrstn_wdma7),
        .o_mclk_y2r_dma                  (mvp_crm_o_mclk_y2r_dma),
        .o_mrstn_y2r_dma                 (mvp_crm_o_mrstn_y2r_dma),
        .o_clk_riscv                     (mvp_crm_o_clk_riscv),
        .o_rstn_riscv                    (mvp_crm_o_rstn_riscv),
        .o_mclk_rdma                     (mvp_crm_o_mclk_rdma),
        .o_mrstn_rdma                    (mvp_crm_o_mrstn_rdma),
        .o_clk_tg                        (mvp_crm_o_clk_tg),
        .o_rstn_tg                       (mvp_crm_o_rstn_tg),
        .o_clk_yuv2rgb                   (mvp_crm_o_clk_yuv2rgb),
        .o_rstn_yuv2rgb                  (mvp_crm_o_rstn_yuv2rgb),
        .o_clk_dvp0                      (mvp_crm_o_clk_dvp0),
        .o_rstn_dvp0                     (mvp_crm_o_rstn_dvp0),
        .o_clk_dvp1                      (mvp_crm_o_clk_dvp1),
        .o_rstn_dvp1                     (mvp_crm_o_rstn_dvp1),
        .o_clk_dvp2                      (mvp_crm_o_clk_dvp2),
        .o_rstn_dvp2                     (mvp_crm_o_rstn_dvp2),
        .o_clk_dvp3                      (mvp_crm_o_clk_dvp3),
        .o_rstn_dvp3                     (mvp_crm_o_rstn_dvp3),
        .o_clk_dvp4                      (mvp_crm_o_clk_dvp4),
        .o_rstn_dvp4                     (mvp_crm_o_rstn_dvp4),
        .o_clk_dvp5                      (mvp_crm_o_clk_dvp5),
        .o_rstn_dvp5                     (mvp_crm_o_rstn_dvp5),
        .o_clk_dvp6                      (mvp_crm_o_clk_dvp6),
        .o_rstn_dvp6                     (mvp_crm_o_rstn_dvp6),
        .o_clk_dvp7                      (mvp_crm_o_clk_dvp7),
        .o_rstn_dvp7                     (mvp_crm_o_rstn_dvp7),
        .o_clk_isp0_clk                  (mvp_crm_o_clk_isp0_clk),
        .o_rstn_isp0_clk                 (mvp_crm_o_rstn_isp0_clk),
        .o_clk_isp1_clk                  (mvp_crm_o_clk_isp1_clk),
        .o_rstn_isp1_clk                 (mvp_crm_o_rstn_isp1_clk),
        .o_clk_isp2_clk                  (mvp_crm_o_clk_isp2_clk),
        .o_rstn_isp2_clk                 (mvp_crm_o_rstn_isp2_clk),
        .o_clk_isp3_clk                  (mvp_crm_o_clk_isp3_clk),
        .o_rstn_isp3_clk                 (mvp_crm_o_rstn_isp3_clk),
        .o_clk_isp4_clk                  (mvp_crm_o_clk_isp4_clk),
        .o_rstn_isp4_clk                 (mvp_crm_o_rstn_isp4_clk),
        .o_clk_isp5_clk                  (mvp_crm_o_clk_isp5_clk),
        .o_rstn_isp5_clk                 (mvp_crm_o_rstn_isp5_clk),
        .o_clk_isp6_clk                  (mvp_crm_o_clk_isp6_clk),
        .o_rstn_isp6_clk                 (mvp_crm_o_rstn_isp6_clk),
        .o_clk_isp7_clk                  (mvp_crm_o_clk_isp7_clk),
        .o_rstn_isp7_clk                 (mvp_crm_o_rstn_isp7_clk),
        .i_scan_mode                     (i_crm_test_mode),
        .i_scan_rstn                     (i_test_rstn),
        .i_test_clk100                   (i_test_clk100),
        .i_test_clk24                    (i_test_clk24),
        .i_test_clk300                   (i_test_clk300)
    );

    tmux_sf_pll2551x_ln28lpp_5000 u_pll_tg (
        .i_tmode                         (i_test_mode),
        .i_norm_p                        (mvp_crm_o_pll_tg_norm_p),
        .i_norm_m                        (mvp_crm_o_pll_tg_norm_m),
        .i_norm_s                        (mvp_crm_o_pll_tg_norm_s),
        .i_norm_lock_con_in              (mvp_crm_o_pll_tg_norm_lock_con_in),
        .i_norm_lock_con_out             (mvp_crm_o_pll_tg_norm_lock_con_out),
        .i_norm_lock_con_dly             (mvp_crm_o_pll_tg_norm_lock_con_dly),
        .i_norm_lock_con_rev             (mvp_crm_o_pll_tg_norm_lock_con_rev),
        .i_norm_tst_afc                  (mvp_crm_o_pll_tg_norm_tst_afc),
        .i_norm_icp                      (mvp_crm_o_pll_tg_norm_icp),
        .i_norm_fin                      (mvp_crm_o_clk_phy_ref),
        .i_norm_resetb                   (mvp_crm_o_pll_tg_norm_resetb),
        .i_norm_bypass                   (mvp_crm_o_pll_tg_norm_bypass),
        .i_norm_tst_en                   (mvp_crm_o_pll_tg_norm_tst_en),
        .i_norm_fsel                     (mvp_crm_o_pll_tg_norm_fsel),
        .i_norm_feed_en                  (mvp_crm_o_pll_tg_norm_feed_en),
        .i_norm_lock_en                  (mvp_crm_o_pll_tg_norm_lock_en),
        .i_norm_afcini_sel               (mvp_crm_o_pll_tg_norm_afcini_sel),
        .i_norm_vcoini_en                (mvp_crm_o_pll_tg_norm_vcoini_en),
        .i_norm_fout_mask                (mvp_crm_o_pll_tg_norm_fout_mask),
        .i_norm_pbias_ctrl               (mvp_crm_o_pll_tg_norm_pbias_ctrl),
        .i_norm_pbias_ctrl_en            (mvp_crm_o_pll_tg_norm_pbias_ctrl_en),
        .i_test_p                        (t_tg_pll_p),
        .i_test_m                        (t_tg_pll_m),
        .i_test_s                        (t_tg_pll_s),
        .i_test_lock_con_in              (t_tg_pll_lock_con_in),
        .i_test_lock_con_out             (t_tg_pll_lock_con_out),
        .i_test_lock_con_dly             (t_tg_pll_lock_con_dly),
        .i_test_lock_con_rev             (t_tg_pll_lock_con_rev),
        .i_test_tst_afc                  (t_tg_pll_tst_afc),
        .i_test_icp                      (t_tg_pll_icp),
        .i_test_fin                      (t_tg_pll_fin),
        .i_test_resetb                   (t_tg_pll_resetb),
        .i_test_bypass                   (t_tg_pll_bypass),
        .i_test_tst_en                   (t_tg_pll_tst_en),
        .i_test_fsel                     (t_tg_pll_fsel),
        .i_test_feed_en                  (t_tg_pll_feed_en),
        .i_test_lock_en                  (t_tg_pll_lock_en),
        .i_test_afcini_sel               (t_tg_pll_afcini_sel),
        .i_test_vcoini_en                (t_tg_pll_vcoini_en),
        .i_test_fout_mask                (t_tg_pll_fout_mask),
        .i_test_pbias_ctrl               (t_tg_pll_pbias_ctrl),
        .i_test_pbias_ctrl_en            (t_tg_pll_pbias_ctrl_en),
        .o_feed_out                      (tg_pll_o_feed_out),
        .o_lock                          (tg_pll_o_lock),
        .o_fout                          (tg_pll_o_fout),
        .o_sync_m_clk_out                (tg_pll_o_sync_m_clk_out),
        .o_afc_code                      (tg_pll_o_afc_code)
    );

    tmux_sf_pll2551x_ln28lpp_5000 u_pll_isp0 (
        .i_tmode                         (i_test_mode),
        .i_norm_p                        (mvp_crm_o_pll_isp0_norm_p),
        .i_norm_m                        (mvp_crm_o_pll_isp0_norm_m),
        .i_norm_s                        (mvp_crm_o_pll_isp0_norm_s),
        .i_norm_lock_con_in              (mvp_crm_o_pll_isp0_norm_lock_con_in),
        .i_norm_lock_con_out             (mvp_crm_o_pll_isp0_norm_lock_con_out),
        .i_norm_lock_con_dly             (mvp_crm_o_pll_isp0_norm_lock_con_dly),
        .i_norm_lock_con_rev             (mvp_crm_o_pll_isp0_norm_lock_con_rev),
        .i_norm_tst_afc                  (mvp_crm_o_pll_isp0_norm_tst_afc),
        .i_norm_icp                      (mvp_crm_o_pll_isp0_norm_icp),
        .i_norm_fin                      (mvp_crm_o_clk_phy_ref),
        .i_norm_resetb                   (mvp_crm_o_pll_isp0_norm_resetb),
        .i_norm_bypass                   (mvp_crm_o_pll_isp0_norm_bypass),
        .i_norm_tst_en                   (mvp_crm_o_pll_isp0_norm_tst_en),
        .i_norm_fsel                     (mvp_crm_o_pll_isp0_norm_fsel),
        .i_norm_feed_en                  (mvp_crm_o_pll_isp0_norm_feed_en),
        .i_norm_lock_en                  (mvp_crm_o_pll_isp0_norm_lock_en),
        .i_norm_afcini_sel               (mvp_crm_o_pll_isp0_norm_afcini_sel),
        .i_norm_vcoini_en                (mvp_crm_o_pll_isp0_norm_vcoini_en),
        .i_norm_fout_mask                (mvp_crm_o_pll_isp0_norm_fout_mask),
        .i_norm_pbias_ctrl               (mvp_crm_o_pll_isp0_norm_pbias_ctrl),
        .i_norm_pbias_ctrl_en            (mvp_crm_o_pll_isp0_norm_pbias_ctrl_en),
        .i_test_p                        (t_isp0_pll_p),
        .i_test_m                        (t_isp0_pll_m),
        .i_test_s                        (t_isp0_pll_s),
        .i_test_lock_con_in              (t_isp0_pll_lock_con_in),
        .i_test_lock_con_out             (t_isp0_pll_lock_con_out),
        .i_test_lock_con_dly             (t_isp0_pll_lock_con_dly),
        .i_test_lock_con_rev             (t_isp0_pll_lock_con_rev),
        .i_test_tst_afc                  (t_isp0_pll_tst_afc),
        .i_test_icp                      (t_isp0_pll_icp),
        .i_test_fin                      (t_isp0_pll_fin),
        .i_test_resetb                   (t_isp0_pll_resetb),
        .i_test_bypass                   (t_isp0_pll_bypass),
        .i_test_tst_en                   (t_isp0_pll_tst_en),
        .i_test_fsel                     (t_isp0_pll_fsel),
        .i_test_feed_en                  (t_isp0_pll_feed_en),
        .i_test_lock_en                  (t_isp0_pll_lock_en),
        .i_test_afcini_sel               (t_isp0_pll_afcini_sel),
        .i_test_vcoini_en                (t_isp0_pll_vcoini_en),
        .i_test_fout_mask                (t_isp0_pll_fout_mask),
        .i_test_pbias_ctrl               (t_isp0_pll_pbias_ctrl),
        .i_test_pbias_ctrl_en            (t_isp0_pll_pbias_ctrl_en),
        .o_feed_out                      (isp0_pll_o_feed_out),
        .o_lock                          (isp0_pll_o_lock),
        .o_fout                          (isp0_pll_o_fout),
        .o_sync_m_clk_out                (isp0_pll_o_sync_m_clk_out),
        .o_afc_code                      (isp0_pll_o_afc_code)
    );

    tmux_sf_pll2551x_ln28lpp_5000 u_pll_isp1 (
        .i_tmode                         (i_test_mode),
        .i_norm_p                        (mvp_crm_o_pll_isp1_norm_p),
        .i_norm_m                        (mvp_crm_o_pll_isp1_norm_m),
        .i_norm_s                        (mvp_crm_o_pll_isp1_norm_s),
        .i_norm_lock_con_in              (mvp_crm_o_pll_isp1_norm_lock_con_in),
        .i_norm_lock_con_out             (mvp_crm_o_pll_isp1_norm_lock_con_out),
        .i_norm_lock_con_dly             (mvp_crm_o_pll_isp1_norm_lock_con_dly),
        .i_norm_lock_con_rev             (mvp_crm_o_pll_isp1_norm_lock_con_rev),
        .i_norm_tst_afc                  (mvp_crm_o_pll_isp1_norm_tst_afc),
        .i_norm_icp                      (mvp_crm_o_pll_isp1_norm_icp),
        .i_norm_fin                      (mvp_crm_o_clk_phy_ref),
        .i_norm_resetb                   (mvp_crm_o_pll_isp1_norm_resetb),
        .i_norm_bypass                   (mvp_crm_o_pll_isp1_norm_bypass),
        .i_norm_tst_en                   (mvp_crm_o_pll_isp1_norm_tst_en),
        .i_norm_fsel                     (mvp_crm_o_pll_isp1_norm_fsel),
        .i_norm_feed_en                  (mvp_crm_o_pll_isp1_norm_feed_en),
        .i_norm_lock_en                  (mvp_crm_o_pll_isp1_norm_lock_en),
        .i_norm_afcini_sel               (mvp_crm_o_pll_isp1_norm_afcini_sel),
        .i_norm_vcoini_en                (mvp_crm_o_pll_isp1_norm_vcoini_en),
        .i_norm_fout_mask                (mvp_crm_o_pll_isp1_norm_fout_mask),
        .i_norm_pbias_ctrl               (mvp_crm_o_pll_isp1_norm_pbias_ctrl),
        .i_norm_pbias_ctrl_en            (mvp_crm_o_pll_isp1_norm_pbias_ctrl_en),
        .i_test_p                        (t_isp1_pll_p),
        .i_test_m                        (t_isp1_pll_m),
        .i_test_s                        (t_isp1_pll_s),
        .i_test_lock_con_in              (t_isp1_pll_lock_con_in),
        .i_test_lock_con_out             (t_isp1_pll_lock_con_out),
        .i_test_lock_con_dly             (t_isp1_pll_lock_con_dly),
        .i_test_lock_con_rev             (t_isp1_pll_lock_con_rev),
        .i_test_tst_afc                  (t_isp1_pll_tst_afc),
        .i_test_icp                      (t_isp1_pll_icp),
        .i_test_fin                      (t_isp1_pll_fin),
        .i_test_resetb                   (t_isp1_pll_resetb),
        .i_test_bypass                   (t_isp1_pll_bypass),
        .i_test_tst_en                   (t_isp1_pll_tst_en),
        .i_test_fsel                     (t_isp1_pll_fsel),
        .i_test_feed_en                  (t_isp1_pll_feed_en),
        .i_test_lock_en                  (t_isp1_pll_lock_en),
        .i_test_afcini_sel               (t_isp1_pll_afcini_sel),
        .i_test_vcoini_en                (t_isp1_pll_vcoini_en),
        .i_test_fout_mask                (t_isp1_pll_fout_mask),
        .i_test_pbias_ctrl               (t_isp1_pll_pbias_ctrl),
        .i_test_pbias_ctrl_en            (t_isp1_pll_pbias_ctrl_en),
        .o_feed_out                      (isp1_pll_o_feed_out),
        .o_lock                          (isp1_pll_o_lock),
        .o_fout                          (isp1_pll_o_fout),
        .o_sync_m_clk_out                (isp1_pll_o_sync_m_clk_out),
        .o_afc_code                      (isp1_pll_o_afc_code)
    );

    mvp_sub u_mvp_sub (
        .i_clk_phy_ref                   (mvp_crm_o_clk_phy_ref),
        .i_clk_riscv_timer0              (mvp_crm_o_clk_riscv_timer0),
        .i_rstn_riscv_timer0             (mvp_crm_o_rstn_riscv_timer0),
        .i_clk_riscv_timer1              (mvp_crm_o_clk_riscv_timer1),
        .i_rstn_riscv_timer1             (mvp_crm_o_rstn_riscv_timer1),
        .i_clk_cpu2mvp                   (mvp_crm_o_clk_cpu2mvp),
        .i_rstn_cpu2mvp                  (mvp_crm_o_rstn_cpu2mvp),
        .i_sclk_wdma0                    (mvp_crm_o_sclk_wdma0),
        .i_srstn_wdma0                   (mvp_crm_o_srstn_wdma0),
        .i_sclk_wdma1                    (mvp_crm_o_sclk_wdma1),
        .i_srstn_wdma1                   (mvp_crm_o_srstn_wdma1),
        .i_sclk_wdma2                    (mvp_crm_o_sclk_wdma2),
        .i_srstn_wdma2                   (mvp_crm_o_srstn_wdma2),
        .i_sclk_wdma3                    (mvp_crm_o_sclk_wdma3),
        .i_srstn_wdma3                   (mvp_crm_o_srstn_wdma3),
        .i_sclk_wdma4                    (mvp_crm_o_sclk_wdma4),
        .i_srstn_wdma4                   (mvp_crm_o_srstn_wdma4),
        .i_sclk_wdma5                    (mvp_crm_o_sclk_wdma5),
        .i_srstn_wdma5                   (mvp_crm_o_srstn_wdma5),
        .i_sclk_wdma6                    (mvp_crm_o_sclk_wdma6),
        .i_srstn_wdma6                   (mvp_crm_o_srstn_wdma6),
        .i_sclk_wdma7                    (mvp_crm_o_sclk_wdma7),
        .i_srstn_wdma7                   (mvp_crm_o_srstn_wdma7),
        .i_sclk_rdma                     (mvp_crm_o_sclk_rdma),
        .i_srstn_rdma                    (mvp_crm_o_srstn_rdma),
        .i_sclk_y2r_dma                  (mvp_crm_o_sclk_y2r_dma),
        .i_srstn_y2r_dma                 (mvp_crm_o_srstn_y2r_dma),
        .i_clk_mvp2main                  (mvp_crm_o_clk_mvp2main),
        .i_rstn_mvp2main                 (mvp_crm_o_rstn_mvp2main),
        .i_mclk_wdma0                    (mvp_crm_o_mclk_wdma0),
        .i_mrstn_wdma0                   (mvp_crm_o_mrstn_wdma0),
        .i_mclk_wdma1                    (mvp_crm_o_mclk_wdma1),
        .i_mrstn_wdma1                   (mvp_crm_o_mrstn_wdma1),
        .i_mclk_wdma2                    (mvp_crm_o_mclk_wdma2),
        .i_mrstn_wdma2                   (mvp_crm_o_mrstn_wdma2),
        .i_mclk_wdma3                    (mvp_crm_o_mclk_wdma3),
        .i_mrstn_wdma3                   (mvp_crm_o_mrstn_wdma3),
        .i_mclk_wdma4                    (mvp_crm_o_mclk_wdma4),
        .i_mrstn_wdma4                   (mvp_crm_o_mrstn_wdma4),
        .i_mclk_wdma5                    (mvp_crm_o_mclk_wdma5),
        .i_mrstn_wdma5                   (mvp_crm_o_mrstn_wdma5),
        .i_mclk_wdma6                    (mvp_crm_o_mclk_wdma6),
        .i_mrstn_wdma6                   (mvp_crm_o_mrstn_wdma6),
        .i_mclk_wdma7                    (mvp_crm_o_mclk_wdma7),
        .i_mrstn_wdma7                   (mvp_crm_o_mrstn_wdma7),
        .i_mclk_rdma                     (mvp_crm_o_mclk_rdma),
        .i_mrstn_rdma                    (mvp_crm_o_mrstn_rdma),
        .i_mclk_y2r_dma                  (mvp_crm_o_mclk_y2r_dma),
        .i_mrstn_y2r_dma                 (mvp_crm_o_mrstn_y2r_dma),
        .i_clk_riscv                     (mvp_crm_o_clk_riscv),
        .i_rstn_riscv                    (mvp_crm_o_rstn_riscv),
        .i_clk_tg                        (mvp_crm_o_clk_tg),
        .i_rstn_tg                       (mvp_crm_o_rstn_tg),
        .i_clk_yuv2rgb                   (mvp_crm_o_clk_yuv2rgb),
        .i_rstn_yuv2rgb                  (mvp_crm_o_rstn_yuv2rgb),
        .i_clk_dvp0_y                    (mvp_crm_o_clk_dvp0),
        .i_rstn_dvp0_y                   (mvp_crm_o_rstn_dvp0),
        .i_clk_dvp1_y                    (mvp_crm_o_clk_dvp1),
        .i_rstn_dvp1_y                   (mvp_crm_o_rstn_dvp1),
        .i_clk_dvp2_y                    (mvp_crm_o_clk_dvp2),
        .i_rstn_dvp2_y                   (mvp_crm_o_rstn_dvp2),
        .i_clk_dvp3_y                    (mvp_crm_o_clk_dvp3),
        .i_rstn_dvp3_y                   (mvp_crm_o_rstn_dvp3),
        .i_clk_dvp4_y                    (mvp_crm_o_clk_dvp4),
        .i_rstn_dvp4_y                   (mvp_crm_o_rstn_dvp4),
        .i_clk_dvp5_y                    (mvp_crm_o_clk_dvp5),
        .i_rstn_dvp5_y                   (mvp_crm_o_rstn_dvp5),
        .i_clk_dvp6_y                    (mvp_crm_o_clk_dvp6),
        .i_rstn_dvp6_y                   (mvp_crm_o_rstn_dvp6),
        .i_clk_dvp7_y                    (mvp_crm_o_clk_dvp7),
        .i_rstn_dvp7_y                   (mvp_crm_o_rstn_dvp7),
        .i_clk_isp0                      (mvp_crm_o_clk_isp0_clk),
        .i_rstn_isp0                     (mvp_crm_o_rstn_isp0_clk),
        .i_clk_isp1                      (mvp_crm_o_clk_isp1_clk),
        .i_rstn_isp1                     (mvp_crm_o_rstn_isp1_clk),
        .i_clk_isp2                      (mvp_crm_o_clk_isp2_clk),
        .i_rstn_isp2                     (mvp_crm_o_rstn_isp2_clk),
        .i_clk_isp3                      (mvp_crm_o_clk_isp3_clk),
        .i_rstn_isp3                     (mvp_crm_o_rstn_isp3_clk),
        .i_clk_isp4                      (mvp_crm_o_clk_isp4_clk),
        .i_rstn_isp4                     (mvp_crm_o_rstn_isp4_clk),
        .i_clk_isp5                      (mvp_crm_o_clk_isp5_clk),
        .i_rstn_isp5                     (mvp_crm_o_rstn_isp5_clk),
        .i_clk_isp6                      (mvp_crm_o_clk_isp6_clk),
        .i_rstn_isp6                     (mvp_crm_o_rstn_isp6_clk),
        .i_clk_isp7                      (mvp_crm_o_clk_isp7_clk),
        .i_rstn_isp7                     (mvp_crm_o_rstn_isp7_clk),
        .o_irq_wdma_err_00               (o_irq_wdma_err_00),
        .o_irq_wdma_err_01               (o_irq_wdma_err_01),
        .o_irq_wdma_err_02               (o_irq_wdma_err_02),
        .o_irq_wdma_err_03               (o_irq_wdma_err_03),
        .o_irq_wdma_err_04               (o_irq_wdma_err_04),
        .o_irq_wdma_err_05               (o_irq_wdma_err_05),
        .o_irq_wdma_err_06               (o_irq_wdma_err_06),
        .o_irq_wdma_err_07               (o_irq_wdma_err_07),
        .o_irq_wdma_done_00              (o_irq_wdma_done_00),
        .o_irq_wdma_done_01              (o_irq_wdma_done_01),
        .o_irq_wdma_done_02              (o_irq_wdma_done_02),
        .o_irq_wdma_done_03              (o_irq_wdma_done_03),
        .o_irq_wdma_done_04              (o_irq_wdma_done_04),
        .o_irq_wdma_done_05              (o_irq_wdma_done_05),
        .o_irq_wdma_done_06              (o_irq_wdma_done_06),
        .o_irq_wdma_done_07              (o_irq_wdma_done_07),
        .o_irq_rdma_err                  (o_irq_rdma_err),
        .o_irq_rdma_done                 (o_irq_rdma_done),
        .o_irq_rwdma_err                 (o_irq_rwdma_err),
        .o_irq_gwdma_err                 (o_irq_gwdma_err),
        .o_irq_bwdma_err                 (o_irq_bwdma_err),
        .o_irq_rwdma_done                (o_irq_rwdma_done),
        .o_irq_gwdma_done                (o_irq_gwdma_done),
        .o_irq_bwdma_done                (o_irq_bwdma_done),
        .o_irq_qisp0_0                   (o_irq_qisp0_0),
        .o_irq_qisp0_1                   (o_irq_qisp0_1),
        .o_irq_qisp1_0                   (o_irq_qisp1_0),
        .o_irq_qisp1_1                   (o_irq_qisp1_1),
        .i_psel_cpu2mvp                  (i_psel_cpu2mvp),
        .i_penable_cpu2mvp               (i_penable_cpu2mvp),
        .i_pwrite_cpu2mvp                (i_pwrite_cpu2mvp),
        .i_paddr_cpu2mvp                 (i_paddr_cpu2mvp),
        .i_pwdata_cpu2mvp                (i_pwdata_cpu2mvp),
        .o_pready_cpu2mvp                (o_pready_cpu2mvp),
        .o_prdata_cpu2mvp                (o_prdata_cpu2mvp),
        .o_pslverr_cpu2mvp               (o_pslverr_cpu2mvp),
        .o_awid_rgb2main                 (o_awid_rgb2main),
        .o_awvalid_rgb2main              (o_awvalid_rgb2main),
        .i_awready_rgb2main              (i_awready_rgb2main),
        .o_awaddr_rgb2main               (o_awaddr_rgb2main),
        .o_awprot_rgb2main               (o_awprot_rgb2main),
        .o_awlen_rgb2main                (o_awlen_rgb2main),
        .o_awsize_rgb2main               (o_awsize_rgb2main),
        .o_awburst_rgb2main              (o_awburst_rgb2main),
        .o_awlock_rgb2main               (o_awlock_rgb2main),
        .o_awcache_rgb2main              (o_awcache_rgb2main),
        .o_wvalid_rgb2main               (o_wvalid_rgb2main),
        .i_wready_rgb2main               (i_wready_rgb2main),
        .o_wdata_rgb2main                (o_wdata_rgb2main),
        .o_wstrb_rgb2main                (o_wstrb_rgb2main),
        .o_wlast_rgb2main                (o_wlast_rgb2main),
        .i_bid_rgb2main                  (i_bid_rgb2main),
        .i_bvalid_rgb2main               (i_bvalid_rgb2main),
        .o_bready_rgb2main               (o_bready_rgb2main),
        .i_bresp_rgb2main                (i_bresp_rgb2main),
        .o_arid_rgb2main                 (o_arid_rgb2main),
        .o_arprot_rgb2main               (o_arprot_rgb2main),
        .o_arvalid_rgb2main              (o_arvalid_rgb2main),
        .i_arready_rgb2main              (i_arready_rgb2main),
        .o_araddr_rgb2main               (o_araddr_rgb2main),
        .o_arlen_rgb2main                (o_arlen_rgb2main),
        .o_arsize_rgb2main               (o_arsize_rgb2main),
        .o_arburst_rgb2main              (o_arburst_rgb2main),
        .o_arlock_rgb2main               (o_arlock_rgb2main),
        .o_arcache_rgb2main              (o_arcache_rgb2main),
        .i_rvalid_rgb2main               (i_rvalid_rgb2main),
        .i_rid_rgb2main                  (i_rid_rgb2main),
        .o_rready_rgb2main               (o_rready_rgb2main),
        .i_rdata_rgb2main                (i_rdata_rgb2main),
        .i_rlast_rgb2main                (i_rlast_rgb2main),
        .i_rresp_rgb2main                (i_rresp_rgb2main),
        .o_awid_isp2main_0               (o_awid_isp2main_0),
        .o_awvalid_isp2main_0            (o_awvalid_isp2main_0),
        .i_awready_isp2main_0            (i_awready_isp2main_0),
        .o_awaddr_isp2main_0             (o_awaddr_isp2main_0),
        .o_awprot_isp2main_0             (o_awprot_isp2main_0),
        .o_awlen_isp2main_0              (o_awlen_isp2main_0),
        .o_awsize_isp2main_0             (o_awsize_isp2main_0),
        .o_awburst_isp2main_0            (o_awburst_isp2main_0),
        .o_awlock_isp2main_0             (o_awlock_isp2main_0),
        .o_awcache_isp2main_0            (o_awcache_isp2main_0),
        .o_wvalid_isp2main_0             (o_wvalid_isp2main_0),
        .i_wready_isp2main_0             (i_wready_isp2main_0),
        .o_wdata_isp2main_0              (o_wdata_isp2main_0),
        .o_wstrb_isp2main_0              (o_wstrb_isp2main_0),
        .o_wlast_isp2main_0              (o_wlast_isp2main_0),
        .i_bid_isp2main_0                (i_bid_isp2main_0),
        .i_bvalid_isp2main_0             (i_bvalid_isp2main_0),
        .o_bready_isp2main_0             (o_bready_isp2main_0),
        .i_bresp_isp2main_0              (i_bresp_isp2main_0),
        .o_arid_isp2main_0               (o_arid_isp2main_0),
        .o_arprot_isp2main_0             (o_arprot_isp2main_0),
        .o_arvalid_isp2main_0            (o_arvalid_isp2main_0),
        .i_arready_isp2main_0            (i_arready_isp2main_0),
        .o_araddr_isp2main_0             (o_araddr_isp2main_0),
        .o_arlen_isp2main_0              (o_arlen_isp2main_0),
        .o_arsize_isp2main_0             (o_arsize_isp2main_0),
        .o_arburst_isp2main_0            (o_arburst_isp2main_0),
        .o_arlock_isp2main_0             (o_arlock_isp2main_0),
        .o_arcache_isp2main_0            (o_arcache_isp2main_0),
        .i_rid_isp2main_0                (i_rid_isp2main_0),
        .i_rvalid_isp2main_0             (i_rvalid_isp2main_0),
        .o_rready_isp2main_0             (o_rready_isp2main_0),
        .i_rdata_isp2main_0              (i_rdata_isp2main_0),
        .i_rlast_isp2main_0              (i_rlast_isp2main_0),
        .i_rresp_isp2main_0              (i_rresp_isp2main_0),
        .o_awid_isp2main_1               (o_awid_isp2main_1),
        .o_awvalid_isp2main_1            (o_awvalid_isp2main_1),
        .i_awready_isp2main_1            (i_awready_isp2main_1),
        .o_awaddr_isp2main_1             (o_awaddr_isp2main_1),
        .o_awprot_isp2main_1             (o_awprot_isp2main_1),
        .o_awlen_isp2main_1              (o_awlen_isp2main_1),
        .o_awsize_isp2main_1             (o_awsize_isp2main_1),
        .o_awburst_isp2main_1            (o_awburst_isp2main_1),
        .o_awlock_isp2main_1             (o_awlock_isp2main_1),
        .o_awcache_isp2main_1            (o_awcache_isp2main_1),
        .o_wvalid_isp2main_1             (o_wvalid_isp2main_1),
        .i_wready_isp2main_1             (i_wready_isp2main_1),
        .o_wdata_isp2main_1              (o_wdata_isp2main_1),
        .o_wstrb_isp2main_1              (o_wstrb_isp2main_1),
        .o_wlast_isp2main_1              (o_wlast_isp2main_1),
        .i_bid_isp2main_1                (i_bid_isp2main_1),
        .i_bvalid_isp2main_1             (i_bvalid_isp2main_1),
        .o_bready_isp2main_1             (o_bready_isp2main_1),
        .i_bresp_isp2main_1              (i_bresp_isp2main_1),
        .o_arid_isp2main_1               (o_arid_isp2main_1),
        .o_arprot_isp2main_1             (o_arprot_isp2main_1),
        .o_arvalid_isp2main_1            (o_arvalid_isp2main_1),
        .i_arready_isp2main_1            (i_arready_isp2main_1),
        .o_araddr_isp2main_1             (o_araddr_isp2main_1),
        .o_arlen_isp2main_1              (o_arlen_isp2main_1),
        .o_arsize_isp2main_1             (o_arsize_isp2main_1),
        .o_arburst_isp2main_1            (o_arburst_isp2main_1),
        .o_arlock_isp2main_1             (o_arlock_isp2main_1),
        .o_arcache_isp2main_1            (o_arcache_isp2main_1),
        .i_rid_isp2main_1                (i_rid_isp2main_1),
        .i_rvalid_isp2main_1             (i_rvalid_isp2main_1),
        .o_rready_isp2main_1             (o_rready_isp2main_1),
        .i_rdata_isp2main_1              (i_rdata_isp2main_1),
        .i_rlast_isp2main_1              (i_rlast_isp2main_1),
        .i_rresp_isp2main_1              (i_rresp_isp2main_1),
        .o_mvp_crm_psel                  (mvp_sub_o_mvp_crm_psel),
        .o_mvp_crm_penable               (mvp_sub_o_mvp_crm_penable),
        .o_mvp_crm_pwrite                (mvp_sub_o_mvp_crm_pwrite),
        .o_mvp_crm_paddr                 (mvp_sub_o_mvp_crm_paddr),
        .o_mvp_crm_pwdata                (mvp_sub_o_mvp_crm_pwdata),
        .i_mvp_crm_prdata                (mvp_sub_i_mvp_crm_prdata),
        .i_mvp_crm_pready                (1'h1),
        .i_mvp_crm_pslverr               (1'h0),
        .i_isp0_cis_dvp_v_y              (i_isp0_cis_dvp_v_y),
        .i_isp0_cis_dvp_h_y              (i_isp0_cis_dvp_h_y),
        .i_isp0_cis_dvp_pv_y             (i_isp0_cis_dvp_pv_y),
        .i_isp0_cis_dvp_p_y              (i_isp0_cis_dvp_p_y),
        .i_isp1_cis_dvp_v_y              (i_isp1_cis_dvp_v_y),
        .i_isp1_cis_dvp_h_y              (i_isp1_cis_dvp_h_y),
        .i_isp1_cis_dvp_pv_y             (i_isp1_cis_dvp_pv_y),
        .i_isp1_cis_dvp_p_y              (i_isp1_cis_dvp_p_y),
        .i_isp2_cis_dvp_v_y              (i_isp2_cis_dvp_v_y),
        .i_isp2_cis_dvp_h_y              (i_isp2_cis_dvp_h_y),
        .i_isp2_cis_dvp_pv_y             (i_isp2_cis_dvp_pv_y),
        .i_isp2_cis_dvp_p_y              (i_isp2_cis_dvp_p_y),
        .i_isp3_cis_dvp_v_y              (i_isp3_cis_dvp_v_y),
        .i_isp3_cis_dvp_h_y              (i_isp3_cis_dvp_h_y),
        .i_isp3_cis_dvp_pv_y             (i_isp3_cis_dvp_pv_y),
        .i_isp3_cis_dvp_p_y              (i_isp3_cis_dvp_p_y),
        .i_isp4_cis_dvp_v_y              (i_isp4_cis_dvp_v_y),
        .i_isp4_cis_dvp_h_y              (i_isp4_cis_dvp_h_y),
        .i_isp4_cis_dvp_pv_y             (i_isp4_cis_dvp_pv_y),
        .i_isp4_cis_dvp_p_y              (i_isp4_cis_dvp_p_y),
        .i_isp5_cis_dvp_v_y              (i_isp5_cis_dvp_v_y),
        .i_isp5_cis_dvp_h_y              (i_isp5_cis_dvp_h_y),
        .i_isp5_cis_dvp_pv_y             (i_isp5_cis_dvp_pv_y),
        .i_isp5_cis_dvp_p_y              (i_isp5_cis_dvp_p_y),
        .i_isp6_cis_dvp_v_y              (i_isp6_cis_dvp_v_y),
        .i_isp6_cis_dvp_h_y              (i_isp6_cis_dvp_h_y),
        .i_isp6_cis_dvp_pv_y             (i_isp6_cis_dvp_pv_y),
        .i_isp6_cis_dvp_p_y              (i_isp6_cis_dvp_p_y),
        .i_isp7_cis_dvp_v_y              (i_isp7_cis_dvp_v_y),
        .i_isp7_cis_dvp_h_y              (i_isp7_cis_dvp_h_y),
        .i_isp7_cis_dvp_pv_y             (i_isp7_cis_dvp_pv_y),
        .i_isp7_cis_dvp_p_y              (i_isp7_cis_dvp_p_y),
        .i_test_mode                     (i_test_mode),
        .i_ema                           (i_ema),
        .o_isp0_i2cm_scl_a               (o_isp0_i2cm_scl_a),
        .o_isp0_i2cm_sda_a               (o_isp0_i2cm_sda_a),
        .o_isp0_i2cm_sda_oe              (o_isp0_i2cm_sda_oe),
        .i_isp0_i2cm_sda_y               (i_isp0_i2cm_sda_y),
        .o_isp1_i2cm_scl_a               (o_isp1_i2cm_scl_a),
        .o_isp1_i2cm_sda_a               (o_isp1_i2cm_sda_a),
        .o_isp1_i2cm_sda_oe              (o_isp1_i2cm_sda_oe),
        .i_isp1_i2cm_sda_y               (i_isp1_i2cm_sda_y),
        .o_isp2_i2cm_scl_a               (o_isp2_i2cm_scl_a),
        .o_isp2_i2cm_sda_a               (o_isp2_i2cm_sda_a),
        .o_isp2_i2cm_sda_oe              (o_isp2_i2cm_sda_oe),
        .i_isp2_i2cm_sda_y               (i_isp2_i2cm_sda_y),
        .o_isp3_i2cm_scl_a               (o_isp3_i2cm_scl_a),
        .o_isp3_i2cm_sda_a               (o_isp3_i2cm_sda_a),
        .o_isp3_i2cm_sda_oe              (o_isp3_i2cm_sda_oe),
        .i_isp3_i2cm_sda_y               (i_isp3_i2cm_sda_y),
        .o_isp4_i2cm_scl_a               (o_isp4_i2cm_scl_a),
        .o_isp4_i2cm_sda_a               (o_isp4_i2cm_sda_a),
        .o_isp4_i2cm_sda_oe              (o_isp4_i2cm_sda_oe),
        .i_isp4_i2cm_sda_y               (i_isp4_i2cm_sda_y),
        .o_isp5_i2cm_scl_a               (o_isp5_i2cm_scl_a),
        .o_isp5_i2cm_sda_a               (o_isp5_i2cm_sda_a),
        .o_isp5_i2cm_sda_oe              (o_isp5_i2cm_sda_oe),
        .i_isp5_i2cm_sda_y               (i_isp5_i2cm_sda_y),
        .o_isp6_i2cm_scl_a               (o_isp6_i2cm_scl_a),
        .o_isp6_i2cm_sda_a               (o_isp6_i2cm_sda_a),
        .o_isp6_i2cm_sda_oe              (o_isp6_i2cm_sda_oe),
        .i_isp6_i2cm_sda_y               (i_isp6_i2cm_sda_y),
        .o_isp7_i2cm_scl_a               (o_isp7_i2cm_scl_a),
        .o_isp7_i2cm_sda_a               (o_isp7_i2cm_sda_a),
        .o_isp7_i2cm_sda_oe              (o_isp7_i2cm_sda_oe),
        .i_isp7_i2cm_sda_y               (i_isp7_i2cm_sda_y),
        .i_i2cs_scl_y                    (i_i2cs_scl_y),
        .o_i2cs_sda_a                    (o_i2cs_sda_a),
        .o_i2cs_sda_oe                   (o_i2cs_sda_oe),
        .i_i2cs_sda_y                    (i_i2cs_sda_y),
        .o_isp0_cis_dvp_p_oe             (o_isp0_cis_dvp_p_oe),
        .o_isp1_cis_dvp_p_oe             (o_isp1_cis_dvp_p_oe),
        .o_isp2_cis_dvp_p_oe             (o_isp2_cis_dvp_p_oe),
        .o_isp3_cis_dvp_p_oe             (o_isp3_cis_dvp_p_oe),
        .o_isp4_cis_dvp_p_oe             (o_isp4_cis_dvp_p_oe),
        .o_isp5_cis_dvp_p_oe             (o_isp5_cis_dvp_p_oe),
        .o_isp6_cis_dvp_p_oe             (o_isp6_cis_dvp_p_oe),
        .o_isp7_cis_dvp_p_oe             (o_isp7_cis_dvp_p_oe),
        .o_isp0_cis_dvp_p_a              (o_isp0_cis_dvp_p_a),
        .o_isp1_cis_dvp_p_a              (o_isp1_cis_dvp_p_a),
        .o_isp2_cis_dvp_p_a              (o_isp2_cis_dvp_p_a),
        .o_isp3_cis_dvp_p_a              (o_isp3_cis_dvp_p_a),
        .o_isp4_cis_dvp_p_a              (o_isp4_cis_dvp_p_a),
        .o_isp5_cis_dvp_p_a              (o_isp5_cis_dvp_p_a),
        .o_isp6_cis_dvp_p_a              (o_isp6_cis_dvp_p_a),
        .o_isp7_cis_dvp_p_a              (o_isp7_cis_dvp_p_a),
        .o_tgclk_a                       (o_tgclk_a),
        .o_tg_dvp_v_a                    (o_tg_dvp_v_a),
        .o_tg_dvp_h_a                    (o_tg_dvp_h_a),
        .o_tg_dvp_p_a                    (o_tg_dvp_p_a),
        .MIPI_CLKP_RX0                   (MIPI_CLKP_RX0),
        .MIPI_CLKN_RX0                   (MIPI_CLKN_RX0),
        .MIPI_DP_RX0                     (MIPI_DP_RX0),
        .MIPI_DN_RX0                     (MIPI_DN_RX0),
        .MIPI_CLKP_RX1                   (MIPI_CLKP_RX1),
        .MIPI_CLKN_RX1                   (MIPI_CLKN_RX1),
        .MIPI_DP_RX1                     (MIPI_DP_RX1),
        .MIPI_DN_RX1                     (MIPI_DN_RX1),
        .MIPI_CLKP_RX2                   (MIPI_CLKP_RX2),
        .MIPI_CLKN_RX2                   (MIPI_CLKN_RX2),
        .MIPI_DP_RX2                     (MIPI_DP_RX2),
        .MIPI_DN_RX2                     (MIPI_DN_RX2),
        .MIPI_CLKP_RX3                   (MIPI_CLKP_RX3),
        .MIPI_CLKN_RX3                   (MIPI_CLKN_RX3),
        .MIPI_DP_RX3                     (MIPI_DP_RX3),
        .MIPI_DN_RX3                     (MIPI_DN_RX3),
        .MIPI_CHIP_EN_MR0                (MIPI_CHIP_EN_MR0),
        .MIPI_HS_CKO_RX0                 (MIPI_HS_CKO_RX0),
        .MIPI_HS_DO_RX0                  (MIPI_HS_DO_RX0),
        .MIPI_TEST_VMON_OUT_RX0          (MIPI_TEST_VMON_OUT_RX0),
        .MIPI_CLKP_RX4                   (MIPI_CLKP_RX4),
        .MIPI_CLKN_RX4                   (MIPI_CLKN_RX4),
        .MIPI_DP_RX4                     (MIPI_DP_RX4),
        .MIPI_DN_RX4                     (MIPI_DN_RX4),
        .MIPI_CLKP_RX5                   (MIPI_CLKP_RX5),
        .MIPI_CLKN_RX5                   (MIPI_CLKN_RX5),
        .MIPI_DP_RX5                     (MIPI_DP_RX5),
        .MIPI_DN_RX5                     (MIPI_DN_RX5),
        .MIPI_CLKP_RX6                   (MIPI_CLKP_RX6),
        .MIPI_CLKN_RX6                   (MIPI_CLKN_RX6),
        .MIPI_DP_RX6                     (MIPI_DP_RX6),
        .MIPI_DN_RX6                     (MIPI_DN_RX6),
        .MIPI_CLKP_RX7                   (MIPI_CLKP_RX7),
        .MIPI_CLKN_RX7                   (MIPI_CLKN_RX7),
        .MIPI_DP_RX7                     (MIPI_DP_RX7),
        .MIPI_DN_RX7                     (MIPI_DN_RX7),
        .MIPI_CHIP_EN_MR1                (MIPI_CHIP_EN_MR1),
        .MIPI_HS_CKO_RX4                 (MIPI_HS_CKO_RX4),
        .MIPI_HS_DO_RX4                  (MIPI_HS_DO_RX4),
        .MIPI_TEST_VMON_OUT_RX4          (MIPI_TEST_VMON_OUT_RX4),
        .MIPI_CHIP_EN_TX                 (MIPI_CHIP_EN_TX),
        .MIPI_CLKP_TX                    (MIPI_CLKP_TX),
        .MIPI_CLKN_TX                    (MIPI_CLKN_TX),
        .MIPI_DP_TX                      (MIPI_DP_TX),
        .MIPI_DN_TX                      (MIPI_DN_TX),
        .MIPI_HS_CKO_TX                  (MIPI_HS_CKO_TX),
        .MIPI_HS_DO_TX                   (MIPI_HS_DO_TX),
        .MIPI_TEST_VMON_OUT_TX           (MIPI_TEST_VMON_OUT_TX),
        .MIPI_TEST_CLK_A0                (MIPI_TEST_CLK_A0),
        .o_awuser_isp2main_0             (o_awuser_isp2main_0),
        .o_awuser_isp2main_1             (o_awuser_isp2main_1),
        .o_awuser_rgb2main               (o_awuser_rgb2main),
        .o_aruser_isp2main_0             (o_aruser_isp2main_0),
        .o_aruser_isp2main_1             (o_aruser_isp2main_1),
        .o_aruser_rgb2main               (o_aruser_rgb2main)
    );

endmodule