module master_axi_128 (
    input             i_aclk   ,
    input             i_aresetn,
    output            o_irq    ,
    output [3:0]      o_awid   ,
    output [31:0]     o_awaddr ,
    output [3:0]      o_awlen  ,
    output [2:0]      o_awsize ,
    output [1:0]      o_awburst,
    output [1:0]      o_awlock ,
    output [3:0]      o_awcache,
    output [2:0]      o_awprot ,
    output            o_awvalid,
    input             i_awready,
    output [3:0]      o_wid    ,
    output [127:0]    o_wdata  ,
    output [15:0]     o_wstrb  ,
    output            o_wlast  ,
    output            o_wvalid ,
    input             i_wready ,
    input  [3:0]      i_bid    ,
    input  [1:0]      i_bresp  ,
    input             i_bvalid ,
    output            o_bready ,
    output [3:0]      o_arid   ,
    output [31:0]     o_araddr ,
    output [3:0]      o_arlen  ,
    output [2:0]      o_arsize ,
    output [1:0]      o_arburst,
    output [1:0]      o_arlock ,
    output [3:0]      o_arcache,
    output [2:0]      o_arprot ,
    output            o_arvalid,
    input             i_arready,
    input  [3:0]      i_rid    ,
    input  [127:0]    i_rdata  ,
    input  [1:0]      i_rresp  ,
    input             i_rlast  ,
    input             i_rvalid ,
    output            o_rready 
);


endmodule