module core_top (
    input   [  7:  0]  i_gpio14_y,
    output  [  7:  0]  o_gpio14_a,
    output  [  7:  0]  o_gpio14_oe,
    input   [  7:  0]  i_gpio12_y,
    output  [  7:  0]  o_gpio12_a,
    output  [  7:  0]  o_gpio12_oe,
    input   [  1:  0]  i_boot_sel_y,
    output  [  1:  0]  o_boot_sel_a,
    output  [  1:  0]  o_boot_sel_oe,
    input   [  7:  0]  i_gpio3_y,
    output  [  7:  0]  o_gpio3_a,
    output  [  7:  0]  o_gpio3_oe,
    input   [  7:  0]  i_gpio7_y,
    output  [  7:  0]  o_gpio7_a,
    output  [  7:  0]  o_gpio7_oe,
    input   [  2:  0]  i_boot_cfg_y,
    output  [  2:  0]  o_boot_cfg_a,
    output  [  2:  0]  o_boot_cfg_oe,
    input   [  7:  0]  i_gpio1_y,
    output  [  7:  0]  o_gpio1_a,
    output  [  7:  0]  o_gpio1_oe,
    input   [  7:  0]  i_gpio9_y,
    output  [  7:  0]  o_gpio9_a,
    output  [  7:  0]  o_gpio9_oe,
    input   [  7:  0]  i_gpio15_y,
    output  [  7:  0]  o_gpio15_a,
    output  [  7:  0]  o_gpio15_oe,
    input   [  7:  0]  i_gpio11_y,
    output  [  7:  0]  o_gpio11_a,
    output  [  7:  0]  o_gpio11_oe,
    input   [  7:  0]  i_gpio8_y,
    output  [  7:  0]  o_gpio8_a,
    output  [  7:  0]  o_gpio8_oe,
    input   [  7:  0]  i_gpio4_y,
    output  [  7:  0]  o_gpio4_a,
    output  [  7:  0]  o_gpio4_oe,
    output  [ 15:  0]  o_tracedata_a,
    input   [  7:  0]  i_gpio17_y,
    output  [  7:  0]  o_gpio17_a,
    output  [  7:  0]  o_gpio17_oe,
    input   [  7:  0]  i_gpio13_y,
    output  [  7:  0]  o_gpio13_a,
    output  [  7:  0]  o_gpio13_oe,
    input   [  7:  0]  i_gpio16_y,
    output  [  7:  0]  o_gpio16_a,
    output  [  7:  0]  o_gpio16_oe,
    input   [  7:  0]  i_gpio10_y,
    output  [  7:  0]  o_gpio10_a,
    output  [  7:  0]  o_gpio10_oe,
    input   [  7:  0]  i_gpio2_y,
    output  [  7:  0]  o_gpio2_a,
    output  [  7:  0]  o_gpio2_oe,
    input   [  7:  0]  i_gpio5_y,
    output  [  7:  0]  o_gpio5_a,
    output  [  7:  0]  o_gpio5_oe,
    input   [  7:  0]  i_gpio0_y,
    output  [  7:  0]  o_gpio0_a,
    output  [  7:  0]  o_gpio0_oe,
    input   [  7:  0]  i_gpio6_y,
    output  [  7:  0]  o_gpio6_a,
    output  [  7:  0]  o_gpio6_oe,
    input   [  7:  0]  i_gpio18_y,
    output  [  7:  0]  o_gpio18_a,
    output  [  7:  0]  o_gpio18_oe,
    input   [  7:  0]  i_gpio19_y,
    output  [  7:  0]  o_gpio19_a,
    output  [  7:  0]  o_gpio19_oe,
    input              i_i2c0_scl_y,
    output             o_i2c0_scl_a,
    output             o_i2c0_scl_oe,
    input              i_i2c0_sda_y,
    output             o_i2c0_sda_a,
    output             o_i2c0_sda_oe,
    input              i_i2c1_scl_y,
    output             o_i2c1_scl_a,
    output             o_i2c1_scl_oe,
    input              i_i2c1_sda_y,
    output             o_i2c1_sda_a,
    output             o_i2c1_sda_oe,
    input              i_i2c2_scl_y,
    output             o_i2c2_scl_a,
    output             o_i2c2_scl_oe,
    input              i_i2c2_sda_y,
    output             o_i2c2_sda_a,
    output             o_i2c2_sda_oe,
    input              i_i2c3_scl_y,
    output             o_i2c3_scl_a,
    output             o_i2c3_scl_oe,
    input              i_i2c3_sda_y,
    output             o_i2c3_sda_a,
    output             o_i2c3_sda_oe,
    input              i_i2s0_bck_y,
    output             o_i2s0_bck_a,
    output             o_i2s0_bck_oe,
    input              i_i2s0_codck_y,
    output             o_i2s0_codck_a,
    output             o_i2s0_codck_oe,
    input              i_i2s0_lrck_y,
    output             o_i2s0_lrck_a,
    output             o_i2s0_lrck_oe,
    input              i_i2s0_rx_y,
    output             o_i2s0_tx_a,
    input              i_i2s1_bck_y,
    output             o_i2s1_bck_a,
    output             o_i2s1_bck_oe,
    input              i_i2s1_codck_y,
    output             o_i2s1_codck_a,
    output             o_i2s1_codck_oe,
    input              i_i2s1_lrck_y,
    output             o_i2s1_lrck_a,
    output             o_i2s1_lrck_oe,
    input              i_i2s1_rx_y,
    output             o_i2s1_tx_a,
    input              i_jtag_ntrst_cs_y,
    input              i_jtag_tck_cs_swclk_y,
    input              i_jtag_tdi_cs_y,
    input              i_jtag_tdo_cs_swo_y,
    output             o_jtag_tdo_cs_swo_a,
    output             o_jtag_tdo_cs_swo_oe,
    input              i_jtag_tms_cs_swdio_y,
    output             o_jtag_tms_cs_swdio_a,
    output             o_jtag_tms_cs_swdio_oe,
    input              i_ssp0_clk_y,
    output             o_ssp0_clk_a,
    output             o_ssp0_clk_oe,
    input              i_ssp0_csn_y,
    output             o_ssp0_csn_a,
    output             o_ssp0_csn_oe,
    input              i_ssp0_rx_y,
    output             o_ssp0_tx_a,
    input              i_ssp1_clk_y,
    output             o_ssp1_clk_a,
    output             o_ssp1_clk_oe,
    input              i_ssp1_csn_y,
    output             o_ssp1_csn_a,
    output             o_ssp1_csn_oe,
    input              i_ssp1_rx_y,
    output             o_ssp1_tx_a,
    input              i_ssp2_clk_y,
    output             o_ssp2_clk_a,
    output             o_ssp2_clk_oe,
    input              i_ssp2_csn_y,
    output             o_ssp2_csn_a,
    output             o_ssp2_csn_oe,
    input              i_ssp2_rx_y,
    output             o_ssp2_tx_a,
    input              i_ssp3_clk_y,
    output             o_ssp3_clk_a,
    output             o_ssp3_clk_oe,
    input              i_ssp3_csn_y,
    output             o_ssp3_csn_a,
    output             o_ssp3_csn_oe,
    input              i_ssp3_rx_y,
    output             o_ssp3_tx_a,
    output             o_traceclk_a,
    output             o_tracectl_a,
    input              i_uart0_rxd_y,
    output             o_uart0_txd_a,
    input              i_uart1_rxd_y,
    output             o_uart1_txd_a,
    input              i_uart2_rxd_y,
    output             o_uart2_txd_a,
    input              i_uart3_rxd_y,
    output             o_uart3_txd_a,
    input              rtc_xin_CK,
    input              xin_CK,
    output  [229:  0]  control_DS0,
    output  [229:  0]  control_DS1,
    output  [229:  0]  control_PE,
    output  [229:  0]  control_PS,
    output  [229:  0]  control_IS,
    output  [229:  0]  control_SR,
    output  [460:  0]  func_sel,
    output  [920:  0]  test_sel,
    output  [230:  0]  func_test_sel
);

    wire    [374:0]  NC_in;
    wire    [704:0]  NC_out;


    peri_hpdf u_peri_hpdf (
        .i_gpio14_y             (i_gpio14_y),
        .o_gpio14_a             (o_gpio14_a),
        .o_gpio14_oe            (o_gpio14_oe),
        .i_gpio12_y             (i_gpio12_y),
        .o_gpio12_a             (o_gpio12_a),
        .o_gpio12_oe            (o_gpio12_oe),
        .i_boot_sel_y           (i_boot_sel_y),
        .o_boot_sel_a           (o_boot_sel_a),
        .o_boot_sel_oe          (o_boot_sel_oe),
        .i_gpio3_y              (i_gpio3_y),
        .o_gpio3_a              (o_gpio3_a),
        .o_gpio3_oe             (o_gpio3_oe),
        .i_gpio7_y              (i_gpio7_y),
        .o_gpio7_a              (o_gpio7_a),
        .o_gpio7_oe             (o_gpio7_oe),
        .i_boot_cfg_y           (i_boot_cfg_y),
        .o_boot_cfg_a           (o_boot_cfg_a),
        .o_boot_cfg_oe          (o_boot_cfg_oe),
        .o_irq_imsi             (NC_out[0]),
        .i_gpio1_y              (i_gpio1_y),
        .o_gpio1_a              (o_gpio1_a),
        .o_gpio1_oe             (o_gpio1_oe),
        .i_gpio9_y              (i_gpio9_y),
        .o_gpio9_a              (o_gpio9_a),
        .o_gpio9_oe             (o_gpio9_oe),
        .i_gpio15_y             (i_gpio15_y),
        .o_gpio15_a             (o_gpio15_a),
        .o_gpio15_oe            (o_gpio15_oe),
        .i_gpio11_y             (i_gpio11_y),
        .o_gpio11_a             (o_gpio11_a),
        .o_gpio11_oe            (o_gpio11_oe),
        .i_gpio8_y              (i_gpio8_y),
        .o_gpio8_a              (o_gpio8_a),
        .o_gpio8_oe             (o_gpio8_oe),
        .i_gpio4_y              (i_gpio4_y),
        .o_gpio4_a              (o_gpio4_a),
        .o_gpio4_oe             (o_gpio4_oe),
        .i_aclk                 (NC_in[0]),
        .i_aresetn              (NC_in[1]),
        .i_peri_awid            (NC_in[5:2]),
        .i_peri_awaddr          (NC_in[37:6]),
        .i_peri_awlen           (NC_in[41:38]),
        .i_peri_awsize          (NC_in[44:42]),
        .i_peri_awburst         (NC_in[46:45]),
        .i_peri_awlock          (NC_in[48:47]),
        .i_peri_awcache         (NC_in[52:49]),
        .i_peri_awprot          (NC_in[55:53]),
        .i_peri_awvalid         (NC_in[56]),
        .o_peri_awready         (NC_out[1]),
        .i_peri_wid             (NC_in[60:57]),
        .i_peri_wdata           (NC_in[188:61]),
        .i_peri_wstrb           (NC_in[204:189]),
        .i_peri_wlast           (NC_in[205]),
        .i_peri_wvalid          (NC_in[206]),
        .o_peri_wready          (NC_out[2]),
        .o_peri_bid             (NC_out[6:3]),
        .o_peri_bresp           (NC_out[8:7]),
        .o_peri_bvalid          (NC_out[9]),
        .i_peri_bready          (NC_in[207]),
        .i_peri_arid            (NC_in[211:208]),
        .i_peri_araddr          (NC_in[243:212]),
        .i_peri_arlen           (NC_in[247:244]),
        .i_peri_arsize          (NC_in[250:248]),
        .i_peri_arburst         (NC_in[252:251]),
        .i_peri_arlock          (NC_in[254:253]),
        .i_peri_arcache         (NC_in[258:255]),
        .i_peri_arprot          (NC_in[261:259]),
        .i_peri_arvalid         (NC_in[262]),
        .o_peri_arready         (NC_out[10]),
        .o_peri_rid             (NC_out[14:11]),
        .o_peri_rdata           (NC_out[142:15]),
        .o_peri_rresp           (NC_out[144:143]),
        .o_peri_rlast           (NC_out[145]),
        .o_peri_rvalid          (NC_out[146]),
        .i_peri_rready          (NC_in[263]),
        .i_pclk                 (NC_in[264]),
        .i_presetn              (NC_in[265]),
        .o_irq                  (NC_out[147]),
        .o_psel                 (NC_out[148]),
        .o_penable              (NC_out[149]),
        .o_paddr                (NC_out[181:150]),
        .o_pwrite               (NC_out[182]),
        .o_pwdata               (NC_out[214:183]),
        .o_pprot                (NC_out[217:215]),
        .o_pstrb                (NC_out[221:218]),
        .i_prdata               (NC_in[297:266]),
        .i_pready               (NC_in[298]),
        .i_pslverr              (NC_in[299]),
        .o_irq_wdt              (NC_out[222]),
        .o_irq_pmu              (NC_out[223]),
        .o_irq_otp              (NC_out[224])
    );

    cpu_interrupt u_cpu_interrupt (
        .o_soc_irq              (NC_out[704:225]),
        .i_irq_wdt              (NC_in[300]),
        .i_irq_timer0_0         (NC_in[301]),
        .i_irq_timer0_1         (NC_in[302]),
        .i_irq_timer0_2         (NC_in[303]),
        .i_irq_timer0_3         (NC_in[304]),
        .i_irq_timer0_4         (NC_in[305]),
        .i_irq_timer1_0         (NC_in[306]),
        .i_irq_timer1_1         (NC_in[307]),
        .i_irq_timer1_2         (NC_in[308]),
        .i_irq_timer1_3         (NC_in[309]),
        .i_irq_timer1_4         (NC_in[310]),
        .i_irq_timer2_0         (NC_in[311]),
        .i_irq_timer2_1         (NC_in[312]),
        .i_irq_timer2_2         (NC_in[313]),
        .i_irq_timer2_3         (NC_in[314]),
        .i_irq_timer2_4         (NC_in[315]),
        .i_irq_timer3_0         (NC_in[316]),
        .i_irq_timer3_1         (NC_in[317]),
        .i_irq_timer3_2         (NC_in[318]),
        .i_irq_timer3_3         (NC_in[319]),
        .i_irq_timer3_4         (NC_in[320]),
        .i_irq_uart0            (NC_in[321]),
        .i_irq_uart1            (NC_in[322]),
        .i_irq_uart2            (NC_in[323]),
        .i_irq_uart3            (NC_in[324]),
        .i_irq_i2c0             (NC_in[325]),
        .i_irq_i2c1             (NC_in[326]),
        .i_irq_i2c2             (NC_in[327]),
        .i_irq_i2c3             (NC_in[328]),
        .i_irq_ssp0_tx          (NC_in[329]),
        .i_irq_ssp0_rx          (NC_in[330]),
        .i_irq_ssp1_tx          (NC_in[331]),
        .i_irq_ssp1_rx          (NC_in[332]),
        .i_irq_ssp2_tx          (NC_in[333]),
        .i_irq_ssp2_rx          (NC_in[334]),
        .i_irq_ssp3_tx          (NC_in[335]),
        .i_irq_ssp3_rx          (NC_in[336]),
        .i_irq_gpio0            (NC_in[337]),
        .i_irq_gpio1            (NC_in[338]),
        .i_irq_gpio2            (NC_in[339]),
        .i_irq_gpio3            (NC_in[340]),
        .i_irq_rtc_tic_0        (NC_in[341]),
        .i_irq_rtc_tic_1        (NC_in[342]),
        .i_irq_rtc_alarm        (NC_in[343]),
        .i_irq_dma330_0_0       (NC_in[344]),
        .i_irq_dma330_0_1       (NC_in[345]),
        .i_irq_dma330_0_2       (NC_in[346]),
        .i_irq_dma330_0_3       (NC_in[347]),
        .i_irq_dma330_0_4       (NC_in[348]),
        .i_irq_dma330_0_5       (NC_in[349]),
        .i_irq_dma330_0_6       (NC_in[350]),
        .i_irq_dma330_0_7       (NC_in[351]),
        .i_irq_dma330_1_0       (NC_in[352]),
        .i_irq_dma330_1_1       (NC_in[353]),
        .i_irq_dma330_1_2       (NC_in[354]),
        .i_irq_dma330_1_3       (NC_in[355]),
        .i_irq_dma330_1_4       (NC_in[356]),
        .i_irq_dma330_1_5       (NC_in[357]),
        .i_irq_dma330_1_6       (NC_in[358]),
        .i_irq_dma330_1_7       (NC_in[359]),
        .i_irq_dma330_2_0       (NC_in[360]),
        .i_irq_dma330_2_1       (NC_in[361]),
        .i_irq_dma330_2_2       (NC_in[362]),
        .i_irq_dma330_2_3       (NC_in[363]),
        .i_irq_dma330_2_4       (NC_in[364]),
        .i_irq_dma330_2_5       (NC_in[365]),
        .i_irq_dma330_2_6       (NC_in[366]),
        .i_irq_dma330_2_7       (NC_in[367]),
        .i_irq_dma330_0_abort   (NC_in[368]),
        .i_irq_dma330_1_abort   (NC_in[369]),
        .i_irq_dma330_2_abort   (NC_in[370]),
        .i_irq_cti_0            (NC_in[371]),
        .i_irq_cti_1            (NC_in[372]),
        .i_irq_cti_2            (NC_in[373]),
        .i_irq_cti_3            (NC_in[374])
    );

endmodule