//==============================================================================
//
// Project : PNAI70X
//
// Verilog RTL(Behavioral) model
//
// This confidential and proprietary source code may be used only as authorized
// by a licensing agreement from ALPHAHOLDINGS Limited. The entire notice above
// must be reproduced on all authorized copies and copies may only be made to
// the extent permitted by a licensing agreement from ALPHAHOLDINGS Limited.
//
// COPYRIGHT (C) ALPHAHOLDINGS, inc. 2022
//
//==============================================================================
// File name : peri_hpdf
// Version : v1.0
// Description :
// Simulator : NC Verilog
// Created by : SoC Designer
// Date : 2022-04-08  17:4
//==============================================================================

module peri_hpdf (
    input              i_test_mode,
    output             o_i2sbclko_0,
    input              i_i2slrclki_0,
    output             o_i2slrclko_0,
    output             o_i2scodclko_0,
    output             o_txdreq_0,
    input              i_txdack_0,
    output             o_rxdreq_0,
    input              i_rxdack_0,
    output             o_i2scodclkoen_0,
    output             o_i2sbclkoen_0,
    output             o_i2slrclkoen_0,
    input              i_i2ssdi_0,
    output             o_i2ssdo_0,
    output             o_i2sbclko_1,
    input              i_i2slrclki_1,
    output             o_i2slrclko_1,
    output             o_i2scodclko_1,
    output             o_txdreq_1,
    input              i_txdack_1,
    output             o_rxdreq_1,
    input              i_rxdack_1,
    output             o_i2scodclkoen_1,
    output             o_i2sbclkoen_1,
    output             o_i2slrclkoen_1,
    input              i_i2ssdi_1,
    output             o_i2ssdo_1,
    input              i_sclin_0,
    input              i_sdain_0,
    output             o_sclout_0,
    output             o_sdaout_0,
    output             o_int_i2c_0,
    input              i_sclin_1,
    input              i_sdain_1,
    output             o_sclout_1,
    output             o_sdaout_1,
    output             o_int_i2c_1,
    input              i_sclin_2,
    input              i_sdain_2,
    output             o_sclout_2,
    output             o_sdaout_2,
    output             o_int_i2c_2,
    input              i_sclin_3,
    input              i_sdain_3,
    output             o_sclout_3,
    output             o_sdaout_3,
    output             o_int_i2c_3,
    output             o_uarttxdmasreq_0,
    output             o_uartrxdmasreq_0,
    output             o_uarttxdmabreq_0,
    output             o_uartrxdmabreq_0,
    input              i_uarttxdmaclr_0,
    input              i_uartrxdmaclr_0,
    output             o_uartintr_0,
    input              i_uartrxd_0,
    output             o_uarttxd_0,
    output             o_uarttxdmasreq_1,
    output             o_uartrxdmasreq_1,
    output             o_uarttxdmabreq_1,
    output             o_uartrxdmabreq_1,
    input              i_uarttxdmaclr_1,
    input              i_uartrxdmaclr_1,
    output             o_uartintr_1,
    input              i_uartrxd_1,
    output             o_uarttxd_1,
    output             o_uarttxdmasreq_2,
    output             o_uartrxdmasreq_2,
    output             o_uarttxdmabreq_2,
    output             o_uartrxdmabreq_2,
    input              i_uarttxdmaclr_2,
    input              i_uartrxdmaclr_2,
    output             o_uartintr_2,
    input              i_uartrxd_2,
    output             o_uarttxd_2,
    output             o_uarttxdmasreq_3,
    output             o_uartrxdmasreq_3,
    output             o_uarttxdmabreq_3,
    output             o_uartrxdmabreq_3,
    input              i_uarttxdmaclr_3,
    input              i_uartrxdmaclr_3,
    output             o_uartintr_3,
    input              i_uartrxd_3,
    output             o_uarttxd_3,
    output             o_sspintr_0,
    output             o_ssptxdamsreq_0,
    output             o_ssprxdmasreq_0,
    output             o_ssptxdmabreq_0,
    output             o_ssprxdmabreq_0,
    input              i_ssptxdmaclr_0,
    input              i_ssprxdmaclr_0,
    output             o_sspfssout_0,
    output             o_sspclkout_0,
    input              i_ssprxd_0,
    output             o_ssptxd_0,
    output             o_nsspctloe_0,
    input              i_sspfssin_0,
    input              i_sspclkin_0,
    output             o_nsspoe_0,
    output             o_sspintr_1,
    output             o_ssptxdamsreq_1,
    output             o_ssprxdmasreq_1,
    output             o_ssptxdmabreq_1,
    output             o_ssprxdmabreq_1,
    input              i_ssptxdmaclr_1,
    input              i_ssprxdmaclr_1,
    output             o_sspfssout_1,
    output             o_sspclkout_1,
    input              i_ssprxd_1,
    output             o_ssptxd_1,
    output             o_nsspctloe_1,
    input              i_sspfssin_1,
    input              i_sspclkin_1,
    output             o_nsspoe_10,
    output             o_sspintr_2,
    output             o_ssptxdamsreq_2,
    output             o_ssprxdmasreq_2,
    output             o_ssptxdmabreq_2,
    output             o_ssprxdmabreq_2,
    input              i_ssptxdmaclr_2,
    input              i_ssprxdmaclr_2,
    output             o_sspfssout_2,
    output             o_sspclkout_2,
    input              i_ssprxd_2,
    output             o_ssptxd_2,
    output             o_nsspctloe_2,
    input              i_sspfssin_2,
    input              i_sspclkin_2,
    output             o_nsspoe_2,
    output             o_sspintr_3,
    output             o_ssptxdamsreq_3,
    output             o_ssprxdmasreq_3,
    output             o_ssptxdmabreq_3,
    output             o_ssprxdmabreq_3,
    input              i_ssptxdmaclr_3,
    input              i_ssprxdmaclr_3,
    output             o_sspfssout_3,
    output             o_sspclkout_3,
    input              i_ssprxd_3,
    output             o_ssptxd_3,
    output             o_nsspctloe_3,
    input              i_sspfssin_3,
    input              i_sspclkin_3,
    output             o_nsspoe_3,
    output  [  4:  0]  o_tintr_0,
    output  [  4:  0]  o_tintr_1,
    output  [  4:  0]  o_tintr_2,
    output  [  4:  0]  o_tintr_3,
    output             o_gpiointr_0,
    output  [  7:  0]  o_ngpen_0,
    output  [  7:  0]  o_gpout_0,
    input   [  7:  0]  i_gpin_0,
    output             o_gpiointr_1,
    output  [  7:  0]  o_ngpen_1,
    output  [  7:  0]  o_gpout_1,
    input   [  7:  0]  i_gpin_1,
    output             o_gpiointr_2,
    output  [  7:  0]  o_ngpen_2,
    output  [  7:  0]  o_gpout_2,
    input   [  7:  0]  i_gpin_2,
    output             o_gpiointr_3,
    output  [  7:  0]  o_ngpen_3,
    output  [  7:  0]  o_gpout_3,
    input   [  7:  0]  i_gpin_3,
    output             o_gpiointr_4,
    output  [  7:  0]  o_ngpen_4,
    output  [  7:  0]  o_gpout_4,
    input   [  7:  0]  i_gpin_4,
    output             o_gpiointr_5,
    output  [  7:  0]  o_ngpen_5,
    output  [  7:  0]  o_gpout_5,
    input   [  7:  0]  i_gpin_5,
    output             o_gpiointr_6,
    output  [  7:  0]  o_ngpen_6,
    output  [  7:  0]  o_gpout_6,
    input   [  7:  0]  i_gpin_6,
    output             o_gpiointr_7,
    output  [  7:  0]  o_ngpen_7,
    output  [  7:  0]  o_gpout_7,
    input   [  7:  0]  i_gpin_7,
    output             o_gpiointr_8,
    output  [  7:  0]  o_ngpen_8,
    output  [  7:  0]  o_gpout_8,
    input   [  7:  0]  i_gpin_8,
    output             o_gpiointr_9,
    output  [  7:  0]  o_ngpen_9,
    output  [  7:  0]  o_gpout_9,
    input   [  7:  0]  i_gpin_9,
    output             o_gpiointr_10,
    output  [  7:  0]  o_ngpen_10,
    output  [  7:  0]  o_gpout_10,
    input   [  7:  0]  i_gpin_10,
    output             o_gpiointr_11,
    output  [  7:  0]  o_ngpen_11,
    output  [  7:  0]  o_gpout_11,
    input   [  7:  0]  i_gpin_11,
    output             o_gpiointr_12,
    output  [  7:  0]  o_ngpen_12,
    output  [  7:  0]  o_gpout_12,
    input   [  7:  0]  i_gpin_12,
    output             o_gpiointr_13,
    output  [  7:  0]  o_ngpen_13,
    output  [  7:  0]  o_gpout_13,
    input   [  7:  0]  i_gpin_13,
    output             o_gpiointr_14,
    output  [  7:  0]  o_ngpen_14,
    output  [  7:  0]  o_gpout_14,
    input   [  7:  0]  i_gpin_14,
    output             o_gpiointr_15,
    output  [  7:  0]  o_ngpen_15,
    output  [  7:  0]  o_gpout_15,
    input   [  7:  0]  i_gpin_15,
    output             o_gpiointr_16,
    output  [  7:  0]  o_ngpen_16,
    output  [  7:  0]  o_gpout_16,
    input   [  7:  0]  i_gpin_16,
    output             o_gpiointr_17,
    output  [  7:  0]  o_ngpen_17,
    output  [  7:  0]  o_gpout_17,
    input   [  7:  0]  i_gpin_17,
    output             o_gpiointr_18,
    output  [  7:  0]  o_ngpen_18,
    output  [  7:  0]  o_gpout_18,
    input   [  7:  0]  i_gpin_18,
    output             o_gpiointr_19,
    output  [  7:  0]  o_ngpen_19,
    output  [  7:  0]  o_gpout_19,
    input   [  7:  0]  i_gpin_19,
    output             o_wdtintr,
    output             o_nresetout,
    output             o_rtc_tic_irq_0,
    output             o_rtc_tic_irq_1,
    output             o_rtc_alarm_irq,
    input              i_osc_rtc,
    output             o_osc_rtc,
    output             o_adc_clk,
    output             o_adc_pd,
    output             o_adc_soc,
    output  [  3:  0]  o_adc_sel,
    input              i_adc_eoc,
    input   [ 11:  0]  i_adc_data,
    input              i_clk_peri_hpdf,
    input              i_rstn_peri_hpdf,
    input              i_clk_peri_codec,
    input              i_test_clk,
    output             o_peri_pselx_codec_hpdf_m3,
    output             o_peri_penable_codec_hpdf_m3,
    output  [ 31:  0]  o_peri_paddr_codec_hpdf_m3,
    output             o_peri_pwrite_codec_hpdf_m3,
    output  [ 31:  0]  o_peri_pwdata_codec_hpdf_m3,
    input   [ 31:  0]  i_peri_prdata_codec_hpdf_m3,
    input              i_peri_pready_codec_hpdf_m3,
    input              i_peri_pslverr_codec_hpdf_m3,
    input   [  4:  0]  i_peri2port_wrap_awid_cpu2peri_m0,
    input   [ 31:  0]  i_peri2port_wrap_awaddr_cpu2peri_m0,
    input   [  7:  0]  i_peri2port_wrap_awlen_cpu2peri_m0,
    input   [  2:  0]  i_peri2port_wrap_awsize_cpu2peri_m0,
    input   [  1:  0]  i_peri2port_wrap_awburst_cpu2peri_m0,
    input              i_peri2port_wrap_awlock_cpu2peri_m0,
    input   [  3:  0]  i_peri2port_wrap_awcache_cpu2peri_m0,
    input   [  2:  0]  i_peri2port_wrap_awprot_cpu2peri_m0,
    input              i_peri2port_wrap_awvalid_cpu2peri_m0,
    output             o_peri2port_wrap_awready_cpu2peri_m0,
    input   [  4:  0]  i_peri2port_wrap_arid_cpu2peri_m0,
    input   [ 31:  0]  i_peri2port_wrap_araddr_cpu2peri_m0,
    input   [  7:  0]  i_peri2port_wrap_arlen_cpu2peri_m0,
    input   [  2:  0]  i_peri2port_wrap_arsize_cpu2peri_m0,
    input   [  1:  0]  i_peri2port_wrap_arburst_cpu2peri_m0,
    input              i_peri2port_wrap_arlock_cpu2peri_m0,
    input   [  3:  0]  i_peri2port_wrap_arcache_cpu2peri_m0,
    input   [  2:  0]  i_peri2port_wrap_arprot_cpu2peri_m0,
    input              i_peri2port_wrap_arvalid_cpu2peri_m0,
    output             o_peri2port_wrap_arready_cpu2peri_m0,
    input   [ 31:  0]  i_peri2port_wrap_wdata_cpu2peri_m0,
    input   [  3:  0]  i_peri2port_wrap_wstrb_cpu2peri_m0,
    input              i_peri2port_wrap_wlast_cpu2peri_m0,
    input              i_peri2port_wrap_wvalid_cpu2peri_m0,
    output             o_peri2port_wrap_wready_cpu2peri_m0,
    output  [  4:  0]  o_peri2port_wrap_bid_cpu2peri_m0,
    output  [  1:  0]  o_peri2port_wrap_bresp_cpu2peri_m0,
    output             o_peri2port_wrap_bvalid_cpu2peri_m0,
    input              i_peri2port_wrap_bready_cpu2peri_m0,
    output  [  4:  0]  o_peri2port_wrap_rid_cpu2peri_m0,
    output  [  1:  0]  o_peri2port_wrap_rresp_cpu2peri_m0,
    output  [ 31:  0]  o_peri2port_wrap_rdata_cpu2peri_m0,
    output             o_peri2port_wrap_rlast_cpu2peri_m0,
    output             o_peri2port_wrap_rvalid_cpu2peri_m0,
    input              i_peri2port_wrap_rready_cpu2peri_m0,
    output             o_peri_pselx_ddr_hpdf_m6,
    output             o_peri_penable_ddr_hpdf_m6,
    output  [ 31:  0]  o_peri_paddr_ddr_hpdf_m6,
    output             o_peri_pwrite_ddr_hpdf_m6,
    output  [ 31:  0]  o_peri_pwdata_ddr_hpdf_m6,
    input   [ 31:  0]  i_peri_prdata_ddr_hpdf_m6,
    input              i_peri_pready_ddr_hpdf_m6,
    input              i_peri_pslverr_ddr_hpdf_m6,
    output             o_peri_pselx_disp_hpdf_m5,
    output             o_peri_penable_disp_hpdf_m5,
    output  [ 31:  0]  o_peri_paddr_disp_hpdf_m5,
    output             o_peri_pwrite_disp_hpdf_m5,
    output  [ 31:  0]  o_peri_pwdata_disp_hpdf_m5,
    input   [ 31:  0]  i_peri_prdata_disp_hpdf_m5,
    input              i_peri_pready_disp_hpdf_m5,
    input              i_peri_pslverr_disp_hpdf_m5,
    output             o_peri_pselx_hsp_hpdf_m2,
    output             o_peri_penable_hsp_hpdf_m2,
    output  [ 31:  0]  o_peri_paddr_hsp_hpdf_m2,
    output             o_peri_pwrite_hsp_hpdf_m2,
    output  [ 31:  0]  o_peri_pwdata_hsp_hpdf_m2,
    input   [ 31:  0]  i_peri_prdata_hsp_hpdf_m2,
    input              i_peri_pready_hsp_hpdf_m2,
    input              i_peri_pslverr_hsp_hpdf_m2,
    output             o_peri_pselx_npu_hpdf_m4,
    output             o_peri_penable_npu_hpdf_m4,
    output  [ 31:  0]  o_peri_paddr_npu_hpdf_m4,
    output             o_peri_pwrite_npu_hpdf_m4,
    output  [ 31:  0]  o_peri_pwdata_npu_hpdf_m4,
    input   [ 31:  0]  i_peri_prdata_npu_hpdf_m4,
    input              i_peri_pready_npu_hpdf_m4,
    input              i_peri_pslverr_npu_hpdf_m4
);

    wire    [31:0]  peri_paddr_peri0_m0;
    wire            peri_pselx_peri0_m0;
    wire            peri_penable_peri0_m0;
    wire            peri_pwrite_peri0_m0;
    wire    [31:0]  peri_prdata_peri0_m0;
    wire    [31:0]  peri_pwdata_peri0_m0;
    wire            peri_pready_peri0_m0;
    wire            peri_pslverr_peri0_m0;
    wire            peri_sub_o_apb_psel;
    wire            peri_sub_o_apb_penable;
    wire            peri_sub_o_apb_pwrite;
    wire    [11:0]  peri_sub_o_apb_paddr;
    wire    [31:0]  peri_sub_o_apb_pwdata;
    wire    [31:0]  peri_sub_i_apb_prdata;
    wire            crm_peri_o_clk_pclk_i2s0;
    wire            crm_peri_o_rstn_u_crg_pclk_i2s0;
    wire            crm_peri_o_clk_pclk_i2s1;
    wire            crm_peri_o_rstn_u_crg_pclk_i2s1;
    wire            crm_peri_o_clk_pclk_i2c0;
    wire            crm_peri_o_rstn_u_crg_pclk_i2c0;
    wire            crm_peri_o_clk_pclk_i2c1;
    wire            crm_peri_o_rstn_u_crg_pclk_i2c1;
    wire            crm_peri_o_clk_pclk_i2c2;
    wire            crm_peri_o_rstn_u_crg_pclk_i2c2;
    wire            crm_peri_o_clk_pclk_i2c3;
    wire            crm_peri_o_rstn_u_crg_pclk_i2c3;
    wire            crm_peri_o_clk_pclk_uart0;
    wire            crm_peri_o_rstn_u_crg_pclk_uart0;
    wire            crm_peri_o_clk_pclk_uart1;
    wire            crm_peri_o_rstn_u_crg_pclk_uart1;
    wire            crm_peri_o_clk_pclk_uart2;
    wire            crm_peri_o_rstn_u_crg_pclk_uart2;
    wire            crm_peri_o_clk_pclk_uart3;
    wire            crm_peri_o_rstn_u_crg_pclk_uart3;
    wire            crm_peri_o_clk_pclk_spi0;
    wire            crm_peri_o_rstn_u_crg_pclk_spi0;
    wire            crm_peri_o_clk_pclk_spi1;
    wire            crm_peri_o_rstn_u_crg_pclk_spi1;
    wire            crm_peri_o_clk_pclk_spi2;
    wire            crm_peri_o_rstn_u_crg_pclk_spi2;
    wire            crm_peri_o_clk_pclk_spi3;
    wire            crm_peri_o_rstn_u_crg_pclk_spi3;
    wire            crm_peri_o_clk_pclk_timer0;
    wire            crm_peri_o_rstn_u_crg_pclk_timer0;
    wire            crm_peri_o_clk_pclk_timer1;
    wire            crm_peri_o_rstn_u_crg_pclk_timer1;
    wire            crm_peri_o_clk_pclk_timer2;
    wire            crm_peri_o_rstn_u_crg_pclk_timer2;
    wire            crm_peri_o_clk_pclk_timer3;
    wire            crm_peri_o_rstn_u_crg_pclk_timer3;
    wire            crm_peri_o_clk_pclk_gpio0;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio0;
    wire            crm_peri_o_clk_pclk_gpio1;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio1;
    wire            crm_peri_o_clk_pclk_gpio2;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio2;
    wire            crm_peri_o_clk_pclk_gpio3;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio3;
    wire            crm_peri_o_clk_pclk_gpio4;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio4;
    wire            crm_peri_o_clk_pclk_gpio5;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio5;
    wire            crm_peri_o_clk_pclk_gpio6;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio6;
    wire            crm_peri_o_clk_pclk_gpio7;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio7;
    wire            crm_peri_o_clk_pclk_gpio8;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio8;
    wire            crm_peri_o_clk_pclk_gpio9;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio9;
    wire            crm_peri_o_clk_pclk_gpio10;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio10;
    wire            crm_peri_o_clk_pclk_gpio11;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio11;
    wire            crm_peri_o_clk_pclk_gpio12;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio12;
    wire            crm_peri_o_clk_pclk_gpio13;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio13;
    wire            crm_peri_o_clk_pclk_gpio14;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio14;
    wire            crm_peri_o_clk_pclk_gpio15;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio15;
    wire            crm_peri_o_clk_pclk_gpio16;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio16;
    wire            crm_peri_o_clk_pclk_gpio17;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio17;
    wire            crm_peri_o_clk_pclk_gpio18;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio18;
    wire            crm_peri_o_clk_pclk_gpio19;
    wire            crm_peri_o_rstn_u_crg_pclk_gpio19;
    wire            crm_peri_o_clk_pclk_wdt;
    wire            crm_peri_o_rstn_u_crg_pclk_wdt;
    wire            crm_peri_o_clk_pclk_rtc;
    wire            crm_peri_o_rstn_u_crg_pclk_rtc;
    wire            crm_peri_o_clk_pclk_adc;
    wire            crm_peri_o_rstn_u_crg_pclk_adc;
    wire            crm_peri_o_clk_peri_bus;
    wire            crm_peri_o_rstn_u_crg_peri_bus;
    wire            crm_peri_o_clk_codec_clk0;
    wire            crm_peri_o_clk_codec_clk1;


    nic400_peri_bus_r0p00 u_peri_bus (
        .paddr_codec_hpdf_m3        (o_peri_paddr_codec_hpdf_m3),
        .pselx_codec_hpdf_m3        (o_peri_pselx_codec_hpdf_m3),
        .penable_codec_hpdf_m3      (o_peri_penable_codec_hpdf_m3),
        .pwrite_codec_hpdf_m3       (o_peri_pwrite_codec_hpdf_m3),
        .prdata_codec_hpdf_m3       (i_peri_prdata_codec_hpdf_m3),
        .pwdata_codec_hpdf_m3       (o_peri_pwdata_codec_hpdf_m3),
        .pready_codec_hpdf_m3       (i_peri_pready_codec_hpdf_m3),
        .pslverr_codec_hpdf_m3      (i_peri_pslverr_codec_hpdf_m3),
        .awid_cpu2peri_s0           (i_peri2port_wrap_awid_cpu2peri_m0),
        .awaddr_cpu2peri_s0         (i_peri2port_wrap_awaddr_cpu2peri_m0),
        .awlen_cpu2peri_s0          (i_peri2port_wrap_awlen_cpu2peri_m0),
        .awsize_cpu2peri_s0         (i_peri2port_wrap_awsize_cpu2peri_m0),
        .awburst_cpu2peri_s0        (i_peri2port_wrap_awburst_cpu2peri_m0),
        .awlock_cpu2peri_s0         (i_peri2port_wrap_awlock_cpu2peri_m0),
        .awcache_cpu2peri_s0        (i_peri2port_wrap_awcache_cpu2peri_m0),
        .awprot_cpu2peri_s0         (i_peri2port_wrap_awprot_cpu2peri_m0),
        .awvalid_cpu2peri_s0        (i_peri2port_wrap_awvalid_cpu2peri_m0),
        .awready_cpu2peri_s0        (o_peri2port_wrap_awready_cpu2peri_m0),
        .wdata_cpu2peri_s0          (i_peri2port_wrap_wdata_cpu2peri_m0),
        .wstrb_cpu2peri_s0          (i_peri2port_wrap_wstrb_cpu2peri_m0),
        .wlast_cpu2peri_s0          (i_peri2port_wrap_wlast_cpu2peri_m0),
        .wvalid_cpu2peri_s0         (i_peri2port_wrap_wvalid_cpu2peri_m0),
        .wready_cpu2peri_s0         (o_peri2port_wrap_wready_cpu2peri_m0),
        .bid_cpu2peri_s0            (o_peri2port_wrap_bid_cpu2peri_m0),
        .bresp_cpu2peri_s0          (o_peri2port_wrap_bresp_cpu2peri_m0),
        .bvalid_cpu2peri_s0         (o_peri2port_wrap_bvalid_cpu2peri_m0),
        .bready_cpu2peri_s0         (i_peri2port_wrap_bready_cpu2peri_m0),
        .arid_cpu2peri_s0           (i_peri2port_wrap_arid_cpu2peri_m0),
        .araddr_cpu2peri_s0         (i_peri2port_wrap_araddr_cpu2peri_m0),
        .arlen_cpu2peri_s0          (i_peri2port_wrap_arlen_cpu2peri_m0),
        .arsize_cpu2peri_s0         (i_peri2port_wrap_arsize_cpu2peri_m0),
        .arburst_cpu2peri_s0        (i_peri2port_wrap_arburst_cpu2peri_m0),
        .arlock_cpu2peri_s0         (i_peri2port_wrap_arlock_cpu2peri_m0),
        .arcache_cpu2peri_s0        (i_peri2port_wrap_arcache_cpu2peri_m0),
        .arprot_cpu2peri_s0         (i_peri2port_wrap_arprot_cpu2peri_m0),
        .arvalid_cpu2peri_s0        (i_peri2port_wrap_arvalid_cpu2peri_m0),
        .arready_cpu2peri_s0        (o_peri2port_wrap_arready_cpu2peri_m0),
        .rid_cpu2peri_s0            (o_peri2port_wrap_rid_cpu2peri_m0),
        .rdata_cpu2peri_s0          (o_peri2port_wrap_rdata_cpu2peri_m0),
        .rresp_cpu2peri_s0          (o_peri2port_wrap_rresp_cpu2peri_m0),
        .rlast_cpu2peri_s0          (o_peri2port_wrap_rlast_cpu2peri_m0),
        .rvalid_cpu2peri_s0         (o_peri2port_wrap_rvalid_cpu2peri_m0),
        .rready_cpu2peri_s0         (i_peri2port_wrap_rready_cpu2peri_m0),
        .paddr_ddr_hpdf_m6          (o_peri_paddr_ddr_hpdf_m6),
        .pselx_ddr_hpdf_m6          (o_peri_pselx_ddr_hpdf_m6),
        .penable_ddr_hpdf_m6        (o_peri_penable_ddr_hpdf_m6),
        .pwrite_ddr_hpdf_m6         (o_peri_pwrite_ddr_hpdf_m6),
        .prdata_ddr_hpdf_m6         (i_peri_prdata_ddr_hpdf_m6),
        .pwdata_ddr_hpdf_m6         (o_peri_pwdata_ddr_hpdf_m6),
        .pready_ddr_hpdf_m6         (i_peri_pready_ddr_hpdf_m6),
        .pslverr_ddr_hpdf_m6        (i_peri_pslverr_ddr_hpdf_m6),
        .paddr_disp_hpdf_m5         (o_peri_paddr_disp_hpdf_m5),
        .pselx_disp_hpdf_m5         (o_peri_pselx_disp_hpdf_m5),
        .penable_disp_hpdf_m5       (o_peri_penable_disp_hpdf_m5),
        .pwrite_disp_hpdf_m5        (o_peri_pwrite_disp_hpdf_m5),
        .prdata_disp_hpdf_m5        (i_peri_prdata_disp_hpdf_m5),
        .pwdata_disp_hpdf_m5        (o_peri_pwdata_disp_hpdf_m5),
        .pready_disp_hpdf_m5        (i_peri_pready_disp_hpdf_m5),
        .pslverr_disp_hpdf_m5       (i_peri_pslverr_disp_hpdf_m5),
        .paddr_hsp_hpdf_m2          (o_peri_paddr_hsp_hpdf_m2),
        .pselx_hsp_hpdf_m2          (o_peri_pselx_hsp_hpdf_m2),
        .penable_hsp_hpdf_m2        (o_peri_penable_hsp_hpdf_m2),
        .pwrite_hsp_hpdf_m2         (o_peri_pwrite_hsp_hpdf_m2),
        .prdata_hsp_hpdf_m2         (i_peri_prdata_hsp_hpdf_m2),
        .pwdata_hsp_hpdf_m2         (o_peri_pwdata_hsp_hpdf_m2),
        .pready_hsp_hpdf_m2         (i_peri_pready_hsp_hpdf_m2),
        .pslverr_hsp_hpdf_m2        (i_peri_pslverr_hsp_hpdf_m2),
        .paddr_npu_hpdf_m4          (o_peri_paddr_npu_hpdf_m4),
        .pselx_npu_hpdf_m4          (o_peri_pselx_npu_hpdf_m4),
        .penable_npu_hpdf_m4        (o_peri_penable_npu_hpdf_m4),
        .pwrite_npu_hpdf_m4         (o_peri_pwrite_npu_hpdf_m4),
        .prdata_npu_hpdf_m4         (i_peri_prdata_npu_hpdf_m4),
        .pwdata_npu_hpdf_m4         (o_peri_pwdata_npu_hpdf_m4),
        .pready_npu_hpdf_m4         (i_peri_pready_npu_hpdf_m4),
        .pslverr_npu_hpdf_m4        (i_peri_pslverr_npu_hpdf_m4),
        .paddr_peri0_m0             (peri_paddr_peri0_m0),
        .pselx_peri0_m0             (peri_pselx_peri0_m0),
        .penable_peri0_m0           (peri_penable_peri0_m0),
        .pwrite_peri0_m0            (peri_pwrite_peri0_m0),
        .prdata_peri0_m0            (peri_prdata_peri0_m0),
        .pwdata_peri0_m0            (peri_pwdata_peri0_m0),
        .pready_peri0_m0            (peri_pready_peri0_m0),
        .pslverr_peri0_m0           (peri_pslverr_peri0_m0),
        .mainclk                    (crm_peri_o_clk_peri_bus),
        .mainclk_r                  (crm_peri_o_clk_peri_bus),
        .mainclken                  (1'h1),
        .mainresetn                 (crm_peri_o_rstn_u_crg_peri_bus),
        .mainresetn_r               (crm_peri_o_rstn_u_crg_peri_bus)
    );

    peri_sub u_peri_sub (
        .i_paddr_peri0_m0           (peri_paddr_peri0_m0),
        .i_pselx_peri0_m0           (peri_pselx_peri0_m0),
        .i_penable_peri0_m0         (peri_penable_peri0_m0),
        .i_pwrite_peri0_m0          (peri_pwrite_peri0_m0),
        .o_prdata_peri0_m0          (peri_prdata_peri0_m0),
        .i_pwdata_peri0_m0          (peri_pwdata_peri0_m0),
        .o_pready_peri0_m0          (peri_pready_peri0_m0),
        .o_pslverr_peri0_m0         (peri_pslverr_peri0_m0),
        .o_apb_psel                 (peri_sub_o_apb_psel),
        .o_apb_penable              (peri_sub_o_apb_penable),
        .o_apb_pwrite               (peri_sub_o_apb_pwrite),
        .o_apb_paddr                (peri_sub_o_apb_paddr),
        .o_apb_pwdata               (peri_sub_o_apb_pwdata),
        .i_apb_prdata               (peri_sub_i_apb_prdata),
        .i_clk_pclk_i2s0            (crm_peri_o_clk_pclk_i2s0),
        .i_rstn_u_crg_pclk_i2s0     (crm_peri_o_rstn_u_crg_pclk_i2s0),
        .i_clk_pclk_i2s1            (crm_peri_o_clk_pclk_i2s1),
        .i_rstn_u_crg_pclk_i2s1     (crm_peri_o_rstn_u_crg_pclk_i2s1),
        .i_clk_pclk_i2c0            (crm_peri_o_clk_pclk_i2c0),
        .i_rstn_u_crg_pclk_i2c0     (crm_peri_o_rstn_u_crg_pclk_i2c0),
        .i_clk_pclk_i2c1            (crm_peri_o_clk_pclk_i2c1),
        .i_rstn_u_crg_pclk_i2c1     (crm_peri_o_rstn_u_crg_pclk_i2c1),
        .i_clk_pclk_i2c2            (crm_peri_o_clk_pclk_i2c2),
        .i_rstn_u_crg_pclk_i2c2     (crm_peri_o_rstn_u_crg_pclk_i2c2),
        .i_clk_pclk_i2c3            (crm_peri_o_clk_pclk_i2c3),
        .i_rstn_u_crg_pclk_i2c3     (crm_peri_o_rstn_u_crg_pclk_i2c3),
        .i_clk_pclk_uart0           (crm_peri_o_clk_pclk_uart0),
        .i_rstn_u_crg_pclk_uart0    (crm_peri_o_rstn_u_crg_pclk_uart0),
        .i_clk_pclk_uart1           (crm_peri_o_clk_pclk_uart1),
        .i_rstn_u_crg_pclk_uart1    (crm_peri_o_rstn_u_crg_pclk_uart1),
        .i_clk_pclk_uart2           (crm_peri_o_clk_pclk_uart2),
        .i_rstn_u_crg_pclk_uart2    (crm_peri_o_rstn_u_crg_pclk_uart2),
        .i_clk_pclk_uart3           (crm_peri_o_clk_pclk_uart3),
        .i_rstn_u_crg_pclk_uart3    (crm_peri_o_rstn_u_crg_pclk_uart3),
        .i_clk_pclk_spi0            (crm_peri_o_clk_pclk_spi0),
        .i_rstn_u_crg_pclk_spi0     (crm_peri_o_rstn_u_crg_pclk_spi0),
        .i_clk_pclk_spi1            (crm_peri_o_clk_pclk_spi1),
        .i_rstn_u_crg_pclk_spi1     (crm_peri_o_rstn_u_crg_pclk_spi1),
        .i_clk_pclk_spi2            (crm_peri_o_clk_pclk_spi2),
        .i_rstn_u_crg_pclk_spi2     (crm_peri_o_rstn_u_crg_pclk_spi2),
        .i_clk_pclk_spi3            (crm_peri_o_clk_pclk_spi3),
        .i_rstn_u_crg_pclk_spi3     (crm_peri_o_rstn_u_crg_pclk_spi3),
        .i_clk_pclk_timer0          (crm_peri_o_clk_pclk_timer0),
        .i_rstn_u_crg_pclk_timer0   (crm_peri_o_rstn_u_crg_pclk_timer0),
        .i_clk_pclk_timer1          (crm_peri_o_clk_pclk_timer1),
        .i_rstn_u_crg_pclk_timer1   (crm_peri_o_rstn_u_crg_pclk_timer1),
        .i_clk_pclk_timer2          (crm_peri_o_clk_pclk_timer2),
        .i_rstn_u_crg_pclk_timer2   (crm_peri_o_rstn_u_crg_pclk_timer2),
        .i_clk_pclk_timer3          (crm_peri_o_clk_pclk_timer3),
        .i_rstn_u_crg_pclk_timer3   (crm_peri_o_rstn_u_crg_pclk_timer3),
        .i_clk_pclk_gpio0           (crm_peri_o_clk_pclk_gpio0),
        .i_rstn_u_crg_pclk_gpio0    (crm_peri_o_rstn_u_crg_pclk_gpio0),
        .i_clk_pclk_gpio1           (crm_peri_o_clk_pclk_gpio1),
        .i_rstn_u_crg_pclk_gpio1    (crm_peri_o_rstn_u_crg_pclk_gpio1),
        .i_clk_pclk_gpio2           (crm_peri_o_clk_pclk_gpio2),
        .i_rstn_u_crg_pclk_gpio2    (crm_peri_o_rstn_u_crg_pclk_gpio2),
        .i_clk_pclk_gpio3           (crm_peri_o_clk_pclk_gpio3),
        .i_rstn_u_crg_pclk_gpio3    (crm_peri_o_rstn_u_crg_pclk_gpio3),
        .i_clk_pclk_gpio4           (crm_peri_o_clk_pclk_gpio4),
        .i_rstn_u_crg_pclk_gpio4    (crm_peri_o_rstn_u_crg_pclk_gpio4),
        .i_clk_pclk_gpio5           (crm_peri_o_clk_pclk_gpio5),
        .i_rstn_u_crg_pclk_gpio5    (crm_peri_o_rstn_u_crg_pclk_gpio5),
        .i_clk_pclk_gpio6           (crm_peri_o_clk_pclk_gpio6),
        .i_rstn_u_crg_pclk_gpio6    (crm_peri_o_rstn_u_crg_pclk_gpio6),
        .i_clk_pclk_gpio7           (crm_peri_o_clk_pclk_gpio7),
        .i_rstn_u_crg_pclk_gpio7    (crm_peri_o_rstn_u_crg_pclk_gpio7),
        .i_clk_pclk_gpio8           (crm_peri_o_clk_pclk_gpio8),
        .i_rstn_u_crg_pclk_gpio8    (crm_peri_o_rstn_u_crg_pclk_gpio8),
        .i_clk_pclk_gpio9           (crm_peri_o_clk_pclk_gpio9),
        .i_rstn_u_crg_pclk_gpio9    (crm_peri_o_rstn_u_crg_pclk_gpio9),
        .i_clk_pclk_gpio10          (crm_peri_o_clk_pclk_gpio10),
        .i_rstn_u_crg_pclk_gpio10   (crm_peri_o_rstn_u_crg_pclk_gpio10),
        .i_clk_pclk_gpio11          (crm_peri_o_clk_pclk_gpio11),
        .i_rstn_u_crg_pclk_gpio11   (crm_peri_o_rstn_u_crg_pclk_gpio11),
        .i_clk_pclk_gpio12          (crm_peri_o_clk_pclk_gpio12),
        .i_rstn_u_crg_pclk_gpio12   (crm_peri_o_rstn_u_crg_pclk_gpio12),
        .i_clk_pclk_gpio13          (crm_peri_o_clk_pclk_gpio13),
        .i_rstn_u_crg_pclk_gpio13   (crm_peri_o_rstn_u_crg_pclk_gpio13),
        .i_clk_pclk_gpio14          (crm_peri_o_clk_pclk_gpio14),
        .i_rstn_u_crg_pclk_gpio14   (crm_peri_o_rstn_u_crg_pclk_gpio14),
        .i_clk_pclk_gpio15          (crm_peri_o_clk_pclk_gpio15),
        .i_rstn_u_crg_pclk_gpio15   (crm_peri_o_rstn_u_crg_pclk_gpio15),
        .i_clk_pclk_gpio16          (crm_peri_o_clk_pclk_gpio16),
        .i_rstn_u_crg_pclk_gpio16   (crm_peri_o_rstn_u_crg_pclk_gpio16),
        .i_clk_pclk_gpio17          (crm_peri_o_clk_pclk_gpio17),
        .i_rstn_u_crg_pclk_gpio17   (crm_peri_o_rstn_u_crg_pclk_gpio17),
        .i_clk_pclk_gpio18          (crm_peri_o_clk_pclk_gpio18),
        .i_rstn_u_crg_pclk_gpio18   (crm_peri_o_rstn_u_crg_pclk_gpio18),
        .i_clk_pclk_gpio19          (crm_peri_o_clk_pclk_gpio19),
        .i_rstn_u_crg_pclk_gpio19   (crm_peri_o_rstn_u_crg_pclk_gpio19),
        .i_clk_pclk_wdt             (crm_peri_o_clk_pclk_wdt),
        .i_rstn_u_crg_pclk_wdt      (crm_peri_o_rstn_u_crg_pclk_wdt),
        .i_clk_pclk_rtc             (crm_peri_o_clk_pclk_rtc),
        .i_rstn_u_crg_pclk_rtc      (crm_peri_o_rstn_u_crg_pclk_rtc),
        .i_clk_pclk_adc             (crm_peri_o_clk_pclk_adc),
        .i_rstn_u_crg_pclk_adc      (crm_peri_o_rstn_u_crg_pclk_adc),
        .i_clk_peri_bus             (crm_peri_o_clk_peri_bus),
        .i_rstn_u_crg_peri_bus      (crm_peri_o_rstn_u_crg_peri_bus),
        .i_scan_tmode               (i_test_mode),
        .o_i2sbclko_0               (o_i2sbclko_0),
        .i_i2slrclki_0              (i_i2slrclki_0),
        .o_i2slrclko_0              (o_i2slrclko_0),
        .i_i2scodclki_0             (crm_peri_o_clk_codec_clk0),
        .o_i2scodclko_0             (o_i2scodclko_0),
        .o_txdreq_0                 (o_txdreq_0),
        .i_txdack_0                 (i_txdack_0),
        .o_rxdreq_0                 (o_rxdreq_0),
        .i_rxdack_0                 (i_rxdack_0),
        .o_i2scodclkoen_0           (o_i2scodclkoen_0),
        .o_i2sbclkoen_0             (o_i2sbclkoen_0),
        .o_i2slrclkoen_0            (o_i2slrclkoen_0),
        .i_i2ssdi_0                 (i_i2ssdi_0),
        .o_i2ssdo_0                 (o_i2ssdo_0),
        .o_i2sbclko_1               (o_i2sbclko_1),
        .i_i2slrclki_1              (i_i2slrclki_1),
        .o_i2slrclko_1              (o_i2slrclko_1),
        .i_i2scodclki_1             (crm_peri_o_clk_codec_clk1),
        .o_i2scodclko_1             (o_i2scodclko_1),
        .o_txdreq_1                 (o_txdreq_1),
        .i_txdack_1                 (i_txdack_1),
        .o_rxdreq_1                 (o_rxdreq_1),
        .i_rxdack_1                 (i_rxdack_1),
        .o_i2scodclkoen_1           (o_i2scodclkoen_1),
        .o_i2sbclkoen_1             (o_i2sbclkoen_1),
        .o_i2slrclkoen_1            (o_i2slrclkoen_1),
        .i_i2ssdi_1                 (i_i2ssdi_1),
        .o_i2ssdo_1                 (o_i2ssdo_1),
        .i_sclin_0                  (i_sclin_0),
        .i_sdain_0                  (i_sdain_0),
        .o_sclout_0                 (o_sclout_0),
        .o_sdaout_0                 (o_sdaout_0),
        .o_int_i2c_0                (o_int_i2c_0),
        .i_sclin_1                  (i_sclin_1),
        .i_sdain_1                  (i_sdain_1),
        .o_sclout_1                 (o_sclout_1),
        .o_sdaout_1                 (o_sdaout_1),
        .o_int_i2c_1                (o_int_i2c_1),
        .i_sclin_2                  (i_sclin_2),
        .i_sdain_2                  (i_sdain_2),
        .o_sclout_2                 (o_sclout_2),
        .o_sdaout_2                 (o_sdaout_2),
        .o_int_i2c_2                (o_int_i2c_2),
        .i_sclin_3                  (i_sclin_3),
        .i_sdain_3                  (i_sdain_3),
        .o_sclout_3                 (o_sclout_3),
        .o_sdaout_3                 (o_sdaout_3),
        .o_int_i2c_3                (o_int_i2c_3),
        .o_uarttxdmasreq_0          (o_uarttxdmasreq_0),
        .o_uartrxdmasreq_0          (o_uartrxdmasreq_0),
        .o_uarttxdmabreq_0          (o_uarttxdmabreq_0),
        .o_uartrxdmabreq_0          (o_uartrxdmabreq_0),
        .i_uarttxdmaclr_0           (i_uarttxdmaclr_0),
        .i_uartrxdmaclr_0           (i_uartrxdmaclr_0),
        .o_uartintr_0               (o_uartintr_0),
        .i_uartrxd_0                (i_uartrxd_0),
        .o_uarttxd_0                (o_uarttxd_0),
        .o_uarttxdmasreq_1          (o_uarttxdmasreq_1),
        .o_uartrxdmasreq_1          (o_uartrxdmasreq_1),
        .o_uarttxdmabreq_1          (o_uarttxdmabreq_1),
        .o_uartrxdmabreq_1          (o_uartrxdmabreq_1),
        .i_uarttxdmaclr_1           (i_uarttxdmaclr_1),
        .i_uartrxdmaclr_1           (i_uartrxdmaclr_1),
        .o_uartintr_1               (o_uartintr_1),
        .i_uartrxd_1                (i_uartrxd_1),
        .o_uarttxd_1                (o_uarttxd_1),
        .o_uarttxdmasreq_2          (o_uarttxdmasreq_2),
        .o_uartrxdmasreq_2          (o_uartrxdmasreq_2),
        .o_uarttxdmabreq_2          (o_uarttxdmabreq_2),
        .o_uartrxdmabreq_2          (o_uartrxdmabreq_2),
        .i_uarttxdmaclr_2           (i_uarttxdmaclr_2),
        .i_uartrxdmaclr_2           (i_uartrxdmaclr_2),
        .o_uartintr_2               (o_uartintr_2),
        .i_uartrxd_2                (i_uartrxd_2),
        .o_uarttxd_2                (o_uarttxd_2),
        .o_uarttxdmasreq_3          (o_uarttxdmasreq_3),
        .o_uartrxdmasreq_3          (o_uartrxdmasreq_3),
        .o_uarttxdmabreq_3          (o_uarttxdmabreq_3),
        .o_uartrxdmabreq_3          (o_uartrxdmabreq_3),
        .i_uarttxdmaclr_3           (i_uarttxdmaclr_3),
        .i_uartrxdmaclr_3           (i_uartrxdmaclr_3),
        .o_uartintr_3               (o_uartintr_3),
        .i_uartrxd_3                (i_uartrxd_3),
        .o_uarttxd_3                (o_uarttxd_3),
        .o_sspintr_0                (o_sspintr_0),
        .o_ssptxdamsreq_0           (o_ssptxdamsreq_0),
        .o_ssprxdmasreq_0           (o_ssprxdmasreq_0),
        .o_ssptxdmabreq_0           (o_ssptxdmabreq_0),
        .o_ssprxdmabreq_0           (o_ssprxdmabreq_0),
        .i_ssptxdmaclr_0            (i_ssptxdmaclr_0),
        .i_ssprxdmaclr_0            (i_ssprxdmaclr_0),
        .o_sspfssout_0              (o_sspfssout_0),
        .o_sspclkout_0              (o_sspclkout_0),
        .i_ssprxd_0                 (i_ssprxd_0),
        .o_ssptxd_0                 (o_ssptxd_0),
        .o_nsspctloe_0              (o_nsspctloe_0),
        .i_sspfssin_0               (i_sspfssin_0),
        .i_sspclkin_0               (i_sspclkin_0),
        .o_nsspoe_0                 (o_nsspoe_0),
        .o_sspintr_1                (o_sspintr_1),
        .o_ssptxdamsreq_1           (o_ssptxdamsreq_1),
        .o_ssprxdmasreq_1           (o_ssprxdmasreq_1),
        .o_ssptxdmabreq_1           (o_ssptxdmabreq_1),
        .o_ssprxdmabreq_1           (o_ssprxdmabreq_1),
        .i_ssptxdmaclr_1            (i_ssptxdmaclr_1),
        .i_ssprxdmaclr_1            (i_ssprxdmaclr_1),
        .o_sspfssout_1              (o_sspfssout_1),
        .o_sspclkout_1              (o_sspclkout_1),
        .i_ssprxd_1                 (i_ssprxd_1),
        .o_ssptxd_1                 (o_ssptxd_1),
        .o_nsspctloe_1              (o_nsspctloe_1),
        .i_sspfssin_1               (i_sspfssin_1),
        .i_sspclkin_1               (i_sspclkin_1),
        .o_nsspoe_10                (o_nsspoe_10),
        .o_sspintr_2                (o_sspintr_2),
        .o_ssptxdamsreq_2           (o_ssptxdamsreq_2),
        .o_ssprxdmasreq_2           (o_ssprxdmasreq_2),
        .o_ssptxdmabreq_2           (o_ssptxdmabreq_2),
        .o_ssprxdmabreq_2           (o_ssprxdmabreq_2),
        .i_ssptxdmaclr_2            (i_ssptxdmaclr_2),
        .i_ssprxdmaclr_2            (i_ssprxdmaclr_2),
        .o_sspfssout_2              (o_sspfssout_2),
        .o_sspclkout_2              (o_sspclkout_2),
        .i_ssprxd_2                 (i_ssprxd_2),
        .o_ssptxd_2                 (o_ssptxd_2),
        .o_nsspctloe_2              (o_nsspctloe_2),
        .i_sspfssin_2               (i_sspfssin_2),
        .i_sspclkin_2               (i_sspclkin_2),
        .o_nsspoe_2                 (o_nsspoe_2),
        .o_sspintr_3                (o_sspintr_3),
        .o_ssptxdamsreq_3           (o_ssptxdamsreq_3),
        .o_ssprxdmasreq_3           (o_ssprxdmasreq_3),
        .o_ssptxdmabreq_3           (o_ssptxdmabreq_3),
        .o_ssprxdmabreq_3           (o_ssprxdmabreq_3),
        .i_ssptxdmaclr_3            (i_ssptxdmaclr_3),
        .i_ssprxdmaclr_3            (i_ssprxdmaclr_3),
        .o_sspfssout_3              (o_sspfssout_3),
        .o_sspclkout_3              (o_sspclkout_3),
        .i_ssprxd_3                 (i_ssprxd_3),
        .o_ssptxd_3                 (o_ssptxd_3),
        .o_nsspctloe_3              (o_nsspctloe_3),
        .i_sspfssin_3               (i_sspfssin_3),
        .i_sspclkin_3               (i_sspclkin_3),
        .o_nsspoe_3                 (o_nsspoe_3),
        .o_tintr_0                  (o_tintr_0),
        .o_tintr_1                  (o_tintr_1),
        .o_tintr_2                  (o_tintr_2),
        .o_tintr_3                  (o_tintr_3),
        .o_gpiointr_0               (o_gpiointr_0),
        .o_ngpen_0                  (o_ngpen_0),
        .o_gpout_0                  (o_gpout_0),
        .i_gpin_0                   (i_gpin_0),
        .o_gpiointr_1               (o_gpiointr_1),
        .o_ngpen_1                  (o_ngpen_1),
        .o_gpout_1                  (o_gpout_1),
        .i_gpin_1                   (i_gpin_1),
        .o_gpiointr_2               (o_gpiointr_2),
        .o_ngpen_2                  (o_ngpen_2),
        .o_gpout_2                  (o_gpout_2),
        .i_gpin_2                   (i_gpin_2),
        .o_gpiointr_3               (o_gpiointr_3),
        .o_ngpen_3                  (o_ngpen_3),
        .o_gpout_3                  (o_gpout_3),
        .i_gpin_3                   (i_gpin_3),
        .o_gpiointr_4               (o_gpiointr_4),
        .o_ngpen_4                  (o_ngpen_4),
        .o_gpout_4                  (o_gpout_4),
        .i_gpin_4                   (i_gpin_4),
        .o_gpiointr_5               (o_gpiointr_5),
        .o_ngpen_5                  (o_ngpen_5),
        .o_gpout_5                  (o_gpout_5),
        .i_gpin_5                   (i_gpin_5),
        .o_gpiointr_6               (o_gpiointr_6),
        .o_ngpen_6                  (o_ngpen_6),
        .o_gpout_6                  (o_gpout_6),
        .i_gpin_6                   (i_gpin_6),
        .o_gpiointr_7               (o_gpiointr_7),
        .o_ngpen_7                  (o_ngpen_7),
        .o_gpout_7                  (o_gpout_7),
        .i_gpin_7                   (i_gpin_7),
        .o_gpiointr_8               (o_gpiointr_8),
        .o_ngpen_8                  (o_ngpen_8),
        .o_gpout_8                  (o_gpout_8),
        .i_gpin_8                   (i_gpin_8),
        .o_gpiointr_9               (o_gpiointr_9),
        .o_ngpen_9                  (o_ngpen_9),
        .o_gpout_9                  (o_gpout_9),
        .i_gpin_9                   (i_gpin_9),
        .o_gpiointr_10              (o_gpiointr_10),
        .o_ngpen_10                 (o_ngpen_10),
        .o_gpout_10                 (o_gpout_10),
        .i_gpin_10                  (i_gpin_10),
        .o_gpiointr_11              (o_gpiointr_11),
        .o_ngpen_11                 (o_ngpen_11),
        .o_gpout_11                 (o_gpout_11),
        .i_gpin_11                  (i_gpin_11),
        .o_gpiointr_12              (o_gpiointr_12),
        .o_ngpen_12                 (o_ngpen_12),
        .o_gpout_12                 (o_gpout_12),
        .i_gpin_12                  (i_gpin_12),
        .o_gpiointr_13              (o_gpiointr_13),
        .o_ngpen_13                 (o_ngpen_13),
        .o_gpout_13                 (o_gpout_13),
        .i_gpin_13                  (i_gpin_13),
        .o_gpiointr_14              (o_gpiointr_14),
        .o_ngpen_14                 (o_ngpen_14),
        .o_gpout_14                 (o_gpout_14),
        .i_gpin_14                  (i_gpin_14),
        .o_gpiointr_15              (o_gpiointr_15),
        .o_ngpen_15                 (o_ngpen_15),
        .o_gpout_15                 (o_gpout_15),
        .i_gpin_15                  (i_gpin_15),
        .o_gpiointr_16              (o_gpiointr_16),
        .o_ngpen_16                 (o_ngpen_16),
        .o_gpout_16                 (o_gpout_16),
        .i_gpin_16                  (i_gpin_16),
        .o_gpiointr_17              (o_gpiointr_17),
        .o_ngpen_17                 (o_ngpen_17),
        .o_gpout_17                 (o_gpout_17),
        .i_gpin_17                  (i_gpin_17),
        .o_gpiointr_18              (o_gpiointr_18),
        .o_ngpen_18                 (o_ngpen_18),
        .o_gpout_18                 (o_gpout_18),
        .i_gpin_18                  (i_gpin_18),
        .o_gpiointr_19              (o_gpiointr_19),
        .o_ngpen_19                 (o_ngpen_19),
        .o_gpout_19                 (o_gpout_19),
        .i_gpin_19                  (i_gpin_19),
        .o_wdtintr                  (o_wdtintr),
        .o_nresetout                (o_nresetout),
        .o_rtc_tic_irq_0            (o_rtc_tic_irq_0),
        .o_rtc_tic_irq_1            (o_rtc_tic_irq_1),
        .o_rtc_alarm_irq            (o_rtc_alarm_irq),
        .i_osc_rtc                  (i_osc_rtc),
        .o_osc_rtc                  (o_osc_rtc),
        .o_adc_clk                  (o_adc_clk),
        .o_adc_pd                   (o_adc_pd),
        .o_adc_soc                  (o_adc_soc),
        .o_adc_sel                  (o_adc_sel),
        .i_adc_eoc                  (i_adc_eoc),
        .i_adc_data                 (i_adc_data)
    );

    pnai70x_crm_peri u_crm_peri (
        .i_apb_pclk                 (i_clk_peri_hpdf),
        .i_apb_prstn                (i_rstn_peri_hpdf),
        .i_apb_psel                 (peri_sub_o_apb_psel),
        .i_apb_penable              (peri_sub_o_apb_penable),
        .i_apb_pwrite               (peri_sub_o_apb_pwrite),
        .i_apb_paddr                (peri_sub_o_apb_paddr),
        .i_apb_pwdata               (peri_sub_o_apb_pwdata),
        .o_apb_prdata               (peri_sub_i_apb_prdata),
        .i_rstn_peri_hpdf           (i_rstn_peri_hpdf),
        .i_clk_peri_hpdf            (i_clk_peri_hpdf),
        .i_clk_peri_codec           (i_clk_peri_codec),
        .o_clk_pclk_i2s0            (crm_peri_o_clk_pclk_i2s0),
        .o_rstn_u_crg_pclk_i2s0     (crm_peri_o_rstn_u_crg_pclk_i2s0),
        .o_clk_pclk_i2s1            (crm_peri_o_clk_pclk_i2s1),
        .o_rstn_u_crg_pclk_i2s1     (crm_peri_o_rstn_u_crg_pclk_i2s1),
        .o_clk_pclk_i2c0            (crm_peri_o_clk_pclk_i2c0),
        .o_rstn_u_crg_pclk_i2c0     (crm_peri_o_rstn_u_crg_pclk_i2c0),
        .o_clk_pclk_i2c1            (crm_peri_o_clk_pclk_i2c1),
        .o_rstn_u_crg_pclk_i2c1     (crm_peri_o_rstn_u_crg_pclk_i2c1),
        .o_clk_pclk_i2c2            (crm_peri_o_clk_pclk_i2c2),
        .o_rstn_u_crg_pclk_i2c2     (crm_peri_o_rstn_u_crg_pclk_i2c2),
        .o_clk_pclk_i2c3            (crm_peri_o_clk_pclk_i2c3),
        .o_rstn_u_crg_pclk_i2c3     (crm_peri_o_rstn_u_crg_pclk_i2c3),
        .o_clk_pclk_uart0           (crm_peri_o_clk_pclk_uart0),
        .o_rstn_u_crg_pclk_uart0    (crm_peri_o_rstn_u_crg_pclk_uart0),
        .o_clk_pclk_uart1           (crm_peri_o_clk_pclk_uart1),
        .o_rstn_u_crg_pclk_uart1    (crm_peri_o_rstn_u_crg_pclk_uart1),
        .o_clk_pclk_uart2           (crm_peri_o_clk_pclk_uart2),
        .o_rstn_u_crg_pclk_uart2    (crm_peri_o_rstn_u_crg_pclk_uart2),
        .o_clk_pclk_uart3           (crm_peri_o_clk_pclk_uart3),
        .o_rstn_u_crg_pclk_uart3    (crm_peri_o_rstn_u_crg_pclk_uart3),
        .o_clk_pclk_spi0            (crm_peri_o_clk_pclk_spi0),
        .o_rstn_u_crg_pclk_spi0     (crm_peri_o_rstn_u_crg_pclk_spi0),
        .o_clk_pclk_spi1            (crm_peri_o_clk_pclk_spi1),
        .o_rstn_u_crg_pclk_spi1     (crm_peri_o_rstn_u_crg_pclk_spi1),
        .o_clk_pclk_spi2            (crm_peri_o_clk_pclk_spi2),
        .o_rstn_u_crg_pclk_spi2     (crm_peri_o_rstn_u_crg_pclk_spi2),
        .o_clk_pclk_spi3            (crm_peri_o_clk_pclk_spi3),
        .o_rstn_u_crg_pclk_spi3     (crm_peri_o_rstn_u_crg_pclk_spi3),
        .o_clk_pclk_timer0          (crm_peri_o_clk_pclk_timer0),
        .o_rstn_u_crg_pclk_timer0   (crm_peri_o_rstn_u_crg_pclk_timer0),
        .o_clk_pclk_timer1          (crm_peri_o_clk_pclk_timer1),
        .o_rstn_u_crg_pclk_timer1   (crm_peri_o_rstn_u_crg_pclk_timer1),
        .o_clk_pclk_timer2          (crm_peri_o_clk_pclk_timer2),
        .o_rstn_u_crg_pclk_timer2   (crm_peri_o_rstn_u_crg_pclk_timer2),
        .o_clk_pclk_timer3          (crm_peri_o_clk_pclk_timer3),
        .o_rstn_u_crg_pclk_timer3   (crm_peri_o_rstn_u_crg_pclk_timer3),
        .o_clk_pclk_gpio0           (crm_peri_o_clk_pclk_gpio0),
        .o_rstn_u_crg_pclk_gpio0    (crm_peri_o_rstn_u_crg_pclk_gpio0),
        .o_clk_pclk_gpio1           (crm_peri_o_clk_pclk_gpio1),
        .o_rstn_u_crg_pclk_gpio1    (crm_peri_o_rstn_u_crg_pclk_gpio1),
        .o_clk_pclk_gpio2           (crm_peri_o_clk_pclk_gpio2),
        .o_rstn_u_crg_pclk_gpio2    (crm_peri_o_rstn_u_crg_pclk_gpio2),
        .o_clk_pclk_gpio3           (crm_peri_o_clk_pclk_gpio3),
        .o_rstn_u_crg_pclk_gpio3    (crm_peri_o_rstn_u_crg_pclk_gpio3),
        .o_clk_pclk_gpio4           (crm_peri_o_clk_pclk_gpio4),
        .o_rstn_u_crg_pclk_gpio4    (crm_peri_o_rstn_u_crg_pclk_gpio4),
        .o_clk_pclk_gpio5           (crm_peri_o_clk_pclk_gpio5),
        .o_rstn_u_crg_pclk_gpio5    (crm_peri_o_rstn_u_crg_pclk_gpio5),
        .o_clk_pclk_gpio6           (crm_peri_o_clk_pclk_gpio6),
        .o_rstn_u_crg_pclk_gpio6    (crm_peri_o_rstn_u_crg_pclk_gpio6),
        .o_clk_pclk_gpio7           (crm_peri_o_clk_pclk_gpio7),
        .o_rstn_u_crg_pclk_gpio7    (crm_peri_o_rstn_u_crg_pclk_gpio7),
        .o_clk_pclk_gpio8           (crm_peri_o_clk_pclk_gpio8),
        .o_rstn_u_crg_pclk_gpio8    (crm_peri_o_rstn_u_crg_pclk_gpio8),
        .o_clk_pclk_gpio9           (crm_peri_o_clk_pclk_gpio9),
        .o_rstn_u_crg_pclk_gpio9    (crm_peri_o_rstn_u_crg_pclk_gpio9),
        .o_clk_pclk_gpio10          (crm_peri_o_clk_pclk_gpio10),
        .o_rstn_u_crg_pclk_gpio10   (crm_peri_o_rstn_u_crg_pclk_gpio10),
        .o_clk_pclk_gpio11          (crm_peri_o_clk_pclk_gpio11),
        .o_rstn_u_crg_pclk_gpio11   (crm_peri_o_rstn_u_crg_pclk_gpio11),
        .o_clk_pclk_gpio12          (crm_peri_o_clk_pclk_gpio12),
        .o_rstn_u_crg_pclk_gpio12   (crm_peri_o_rstn_u_crg_pclk_gpio12),
        .o_clk_pclk_gpio13          (crm_peri_o_clk_pclk_gpio13),
        .o_rstn_u_crg_pclk_gpio13   (crm_peri_o_rstn_u_crg_pclk_gpio13),
        .o_clk_pclk_gpio14          (crm_peri_o_clk_pclk_gpio14),
        .o_rstn_u_crg_pclk_gpio14   (crm_peri_o_rstn_u_crg_pclk_gpio14),
        .o_clk_pclk_gpio15          (crm_peri_o_clk_pclk_gpio15),
        .o_rstn_u_crg_pclk_gpio15   (crm_peri_o_rstn_u_crg_pclk_gpio15),
        .o_clk_pclk_gpio16          (crm_peri_o_clk_pclk_gpio16),
        .o_rstn_u_crg_pclk_gpio16   (crm_peri_o_rstn_u_crg_pclk_gpio16),
        .o_clk_pclk_gpio17          (crm_peri_o_clk_pclk_gpio17),
        .o_rstn_u_crg_pclk_gpio17   (crm_peri_o_rstn_u_crg_pclk_gpio17),
        .o_clk_pclk_gpio18          (crm_peri_o_clk_pclk_gpio18),
        .o_rstn_u_crg_pclk_gpio18   (crm_peri_o_rstn_u_crg_pclk_gpio18),
        .o_clk_pclk_gpio19          (crm_peri_o_clk_pclk_gpio19),
        .o_rstn_u_crg_pclk_gpio19   (crm_peri_o_rstn_u_crg_pclk_gpio19),
        .o_clk_pclk_wdt             (crm_peri_o_clk_pclk_wdt),
        .o_rstn_u_crg_pclk_wdt      (crm_peri_o_rstn_u_crg_pclk_wdt),
        .o_clk_pclk_rtc             (crm_peri_o_clk_pclk_rtc),
        .o_rstn_u_crg_pclk_rtc      (crm_peri_o_rstn_u_crg_pclk_rtc),
        .o_clk_pclk_adc             (crm_peri_o_clk_pclk_adc),
        .o_rstn_u_crg_pclk_adc      (crm_peri_o_rstn_u_crg_pclk_adc),
        .o_clk_peri_bus             (crm_peri_o_clk_peri_bus),
        .o_rstn_u_crg_peri_bus      (crm_peri_o_rstn_u_crg_peri_bus),
        .o_clk_codec_clk0           (crm_peri_o_clk_codec_clk0),
        .o_clk_codec_clk1           (crm_peri_o_clk_codec_clk1),
        .i_scan_clk                 (i_test_clk),
        .i_scan_mode                (i_test_mode),
        .i_scan_rstn                (1'h0)
    );

endmodule