// ==========================================================
//
// (C) COPYRIGHT 2023 Alpha-Holdings INC. ALL RIGHT RESERVED
//
// User : jhkim
// Time : 2023/12/11/14/18/58
// File : core_top.v
//
// ==========================================================

module core_top (
    output  [  3:  0]  o_cm3_tracedata_a,
    input   [  7:  0]  i_gpio5_y,
    output  [  7:  0]  o_gpio5_a,
    output  [  7:  0]  o_gpio5_oe,
    input   [  7:  0]  i_gpio4_y,
    output  [  7:  0]  o_gpio4_a,
    output  [  7:  0]  o_gpio4_oe,
    input   [  7:  0]  i_gpio6_y,
    output  [  7:  0]  o_gpio6_a,
    output  [  7:  0]  o_gpio6_oe,
    input   [  7:  0]  i_gmac_rxd_y,
    input   [  2:  0]  i_boot_cfg_y,
    output  [  4:  0]  o_timer0_a,
    output  [  4:  0]  o_timer1_a,
    input   [  9:  0]  i_isp6_cis_dvp_p_y,
    output  [  9:  0]  o_isp6_cis_dvp_p_a,
    output  [  9:  0]  o_isp6_cis_dvp_p_oe,
    output  [ 31:  0]  o_tg_dvp_p_a,
    input   [  9:  0]  i_isp5_cis_dvp_p_y,
    output  [  9:  0]  o_isp5_cis_dvp_p_a,
    output  [  9:  0]  o_isp5_cis_dvp_p_oe,
    input   [  1:  0]  i_boot_sel_y,
    input   [  7:  0]  i_nfc_data_y,
    output  [  7:  0]  o_nfc_data_a,
    output  [  7:  0]  o_nfc_data_oe,
    input   [  9:  0]  i_isp3_cis_dvp_p_y,
    output  [  9:  0]  o_isp3_cis_dvp_p_a,
    output  [  9:  0]  o_isp3_cis_dvp_p_oe,
    input   [  7:  0]  i_gpio2_y,
    output  [  7:  0]  o_gpio2_a,
    output  [  7:  0]  o_gpio2_oe,
    input   [  9:  0]  i_isp0_cis_dvp_p_y,
    output  [  9:  0]  o_isp0_cis_dvp_p_a,
    output  [  9:  0]  o_isp0_cis_dvp_p_oe,
    input   [  3:  0]  i_sfmc_data_y,
    output  [  3:  0]  o_sfmc_data_a,
    output  [  3:  0]  o_sfmc_data_oe,
    input   [  9:  0]  i_isp4_cis_dvp_p_y,
    output  [  9:  0]  o_isp4_cis_dvp_p_a,
    output  [  9:  0]  o_isp4_cis_dvp_p_oe,
    output  [  7:  0]  o_gmac_txd_a,
    input   [  9:  0]  i_isp7_cis_dvp_p_y,
    output  [  9:  0]  o_isp7_cis_dvp_p_a,
    output  [  9:  0]  o_isp7_cis_dvp_p_oe,
    input   [  7:  0]  i_gpio1_y,
    output  [  7:  0]  o_gpio1_a,
    output  [  7:  0]  o_gpio1_oe,
    input   [  2:  0]  i_gmac_phy_intf_sel_y,
    input   [  7:  0]  i_gpio7_y,
    output  [  7:  0]  o_gpio7_a,
    output  [  7:  0]  o_gpio7_oe,
    input   [  7:  0]  i_gpio3_y,
    output  [  7:  0]  o_gpio3_a,
    output  [  7:  0]  o_gpio3_oe,
    input   [  9:  0]  i_isp1_cis_dvp_p_y,
    output  [  9:  0]  o_isp1_cis_dvp_p_a,
    output  [  9:  0]  o_isp1_cis_dvp_p_oe,
    input   [  9:  0]  i_isp2_cis_dvp_p_y,
    output  [  9:  0]  o_isp2_cis_dvp_p_a,
    output  [  9:  0]  o_isp2_cis_dvp_p_oe,
    input   [  7:  0]  i_gpio0_y,
    output  [  7:  0]  o_gpio0_a,
    output  [  7:  0]  o_gpio0_oe,
    input              i_clk_dvp0_y,
    input              i_clk_dvp1_y,
    input              i_clk_dvp2_y,
    input              i_clk_dvp3_y,
    input              i_clk_dvp4_y,
    input              i_clk_dvp5_y,
    input              i_clk_dvp6_y,
    input              i_clk_dvp7_y,
    output             o_clk_gmac_rmii_a,
    input              i_clk_gmac_rx_y,
    output             o_clk_gmac_rx_a,
    output             o_clk_gmac_rx_oe,
    input              i_clk_gmac_tx_y,
    output             o_clk_gmac_tx_a,
    output             o_clk_gmac_tx_oe,
    output             o_clk_phy_refclk_a,
    output             o_cm3_traceclk_a,
    input              i_gmac_col_y,
    input              i_gmac_crs_y,
    output             o_gmac_mdc_a,
    input              i_gmac_mdio_y,
    output             o_gmac_mdio_a,
    output             o_gmac_mdio_oe,
    input              i_gmac_rx_dv_y,
    input              i_gmac_rx_er_y,
    output             o_gmac_tx_en_a,
    output             o_gmac_tx_er_a,
    input              i_i2c0_scl_y,
    output             o_i2c0_scl_a,
    output             o_i2c0_scl_oe,
    input              i_i2c0_sda_y,
    output             o_i2c0_sda_a,
    output             o_i2c0_sda_oe,
    input              i_i2c1_scl_y,
    output             o_i2c1_scl_a,
    output             o_i2c1_scl_oe,
    input              i_i2c1_sda_y,
    output             o_i2c1_sda_a,
    output             o_i2c1_sda_oe,
    input              i_i2c2_scl_y,
    output             o_i2c2_scl_a,
    output             o_i2c2_scl_oe,
    input              i_i2c2_sda_y,
    output             o_i2c2_sda_a,
    output             o_i2c2_sda_oe,
    input              i_i2c3_scl_y,
    output             o_i2c3_scl_a,
    output             o_i2c3_scl_oe,
    input              i_i2c3_sda_y,
    output             o_i2c3_sda_a,
    output             o_i2c3_sda_oe,
    input              i_i2c4_scl_y,
    output             o_i2c4_scl_a,
    output             o_i2c4_scl_oe,
    input              i_i2c4_sda_y,
    output             o_i2c4_sda_a,
    output             o_i2c4_sda_oe,
    input              i_i2c5_scl_y,
    output             o_i2c5_scl_a,
    output             o_i2c5_scl_oe,
    input              i_i2c5_sda_y,
    output             o_i2c5_sda_a,
    output             o_i2c5_sda_oe,
    input              i_i2c6_scl_y,
    output             o_i2c6_scl_a,
    output             o_i2c6_scl_oe,
    input              i_i2c6_sda_y,
    output             o_i2c6_sda_a,
    output             o_i2c6_sda_oe,
    input              i_i2c7_scl_y,
    output             o_i2c7_scl_a,
    output             o_i2c7_scl_oe,
    input              i_i2c7_sda_y,
    output             o_i2c7_sda_a,
    output             o_i2c7_sda_oe,
    input              i_i2c8_scl_y,
    output             o_i2c8_scl_a,
    output             o_i2c8_scl_oe,
    input              i_i2c8_sda_y,
    output             o_i2c8_sda_a,
    output             o_i2c8_sda_oe,
    input              i_i2c9_scl_y,
    output             o_i2c9_scl_a,
    output             o_i2c9_scl_oe,
    input              i_i2c9_sda_y,
    output             o_i2c9_sda_a,
    output             o_i2c9_sda_oe,
    input              i_i2cs0_scl_y,
    input              i_i2cs0_sda_y,
    output             o_i2cs0_sda_a,
    output             o_i2cs0_sda_oe,
    input              i_i2cs1_scl_y,
    input              i_i2cs1_sda_y,
    output             o_i2cs1_sda_a,
    output             o_i2cs1_sda_oe,
    input              i_isp0_cis_dvp_h_y,
    output             o_isp0_cis_dvp_h_a,
    output             o_isp0_cis_dvp_h_oe,
    input              i_isp0_cis_dvp_pv_y,
    input              i_isp0_cis_dvp_v_y,
    output             o_isp0_cis_dvp_v_a,
    output             o_isp0_cis_dvp_v_oe,
    input              i_isp0_i2cm_scl_y,
    output             o_isp0_i2cm_scl_a,
    output             o_isp0_i2cm_scl_oe,
    input              i_isp0_i2cm_sda_y,
    output             o_isp0_i2cm_sda_a,
    output             o_isp0_i2cm_sda_oe,
    input              i_isp1_cis_dvp_h_y,
    output             o_isp1_cis_dvp_h_a,
    output             o_isp1_cis_dvp_h_oe,
    input              i_isp1_cis_dvp_pv_y,
    input              i_isp1_cis_dvp_v_y,
    output             o_isp1_cis_dvp_v_a,
    output             o_isp1_cis_dvp_v_oe,
    input              i_isp1_i2cm_scl_y,
    output             o_isp1_i2cm_scl_a,
    output             o_isp1_i2cm_scl_oe,
    input              i_isp1_i2cm_sda_y,
    output             o_isp1_i2cm_sda_a,
    output             o_isp1_i2cm_sda_oe,
    input              i_isp2_cis_dvp_h_y,
    output             o_isp2_cis_dvp_h_a,
    output             o_isp2_cis_dvp_h_oe,
    input              i_isp2_cis_dvp_pv_y,
    input              i_isp2_cis_dvp_v_y,
    output             o_isp2_cis_dvp_v_a,
    output             o_isp2_cis_dvp_v_oe,
    input              i_isp2_i2cm_scl_y,
    output             o_isp2_i2cm_scl_a,
    output             o_isp2_i2cm_scl_oe,
    input              i_isp2_i2cm_sda_y,
    output             o_isp2_i2cm_sda_a,
    output             o_isp2_i2cm_sda_oe,
    input              i_isp3_cis_dvp_h_y,
    output             o_isp3_cis_dvp_h_a,
    output             o_isp3_cis_dvp_h_oe,
    input              i_isp3_cis_dvp_pv_y,
    input              i_isp3_cis_dvp_v_y,
    output             o_isp3_cis_dvp_v_a,
    output             o_isp3_cis_dvp_v_oe,
    input              i_isp3_i2cm_scl_y,
    output             o_isp3_i2cm_scl_a,
    output             o_isp3_i2cm_scl_oe,
    input              i_isp3_i2cm_sda_y,
    output             o_isp3_i2cm_sda_a,
    output             o_isp3_i2cm_sda_oe,
    input              i_isp4_cis_dvp_h_y,
    output             o_isp4_cis_dvp_h_a,
    output             o_isp4_cis_dvp_h_oe,
    input              i_isp4_cis_dvp_pv_y,
    input              i_isp4_cis_dvp_v_y,
    output             o_isp4_cis_dvp_v_a,
    output             o_isp4_cis_dvp_v_oe,
    input              i_isp4_i2cm_scl_y,
    output             o_isp4_i2cm_scl_a,
    output             o_isp4_i2cm_scl_oe,
    input              i_isp4_i2cm_sda_y,
    output             o_isp4_i2cm_sda_a,
    output             o_isp4_i2cm_sda_oe,
    input              i_isp5_cis_dvp_h_y,
    output             o_isp5_cis_dvp_h_a,
    output             o_isp5_cis_dvp_h_oe,
    input              i_isp5_cis_dvp_pv_y,
    input              i_isp5_cis_dvp_v_y,
    output             o_isp5_cis_dvp_v_a,
    output             o_isp5_cis_dvp_v_oe,
    input              i_isp5_i2cm_scl_y,
    output             o_isp5_i2cm_scl_a,
    output             o_isp5_i2cm_scl_oe,
    input              i_isp5_i2cm_sda_y,
    output             o_isp5_i2cm_sda_a,
    output             o_isp5_i2cm_sda_oe,
    input              i_isp6_cis_dvp_h_y,
    output             o_isp6_cis_dvp_h_a,
    output             o_isp6_cis_dvp_h_oe,
    input              i_isp6_cis_dvp_pv_y,
    input              i_isp6_cis_dvp_v_y,
    output             o_isp6_cis_dvp_v_a,
    output             o_isp6_cis_dvp_v_oe,
    input              i_isp6_i2cm_scl_y,
    output             o_isp6_i2cm_scl_a,
    output             o_isp6_i2cm_scl_oe,
    input              i_isp6_i2cm_sda_y,
    output             o_isp6_i2cm_sda_a,
    output             o_isp6_i2cm_sda_oe,
    input              i_isp7_cis_dvp_h_y,
    output             o_isp7_cis_dvp_h_a,
    output             o_isp7_cis_dvp_h_oe,
    input              i_isp7_cis_dvp_pv_y,
    input              i_isp7_cis_dvp_v_y,
    output             o_isp7_cis_dvp_v_a,
    output             o_isp7_cis_dvp_v_oe,
    input              i_isp7_i2cm_scl_y,
    output             o_isp7_i2cm_scl_a,
    output             o_isp7_i2cm_scl_oe,
    input              i_isp7_i2cm_sda_y,
    output             o_isp7_i2cm_sda_a,
    output             o_isp7_i2cm_sda_oe,
    input              i_jtag_ntrst_y,
    input              i_jtag_tck_y,
    input              i_jtag_tdi_y,
    input              i_jtag_tdo_y,
    output             o_jtag_tdo_a,
    output             o_jtag_tdo_oe,
    input              i_jtag_tmms_y,
    output             o_jtag_tmms_a,
    output             o_jtag_tmms_oe,
    input              i_mvp0_uart_rx_y,
    output             o_mvp0_uart_tx_a,
    input              i_mvp1_uart_rx_y,
    output             o_mvp1_uart_tx_a,
    output             o_nfc_ale_a,
    input              i_nfc_cfgaddrcycle_y,
    input              i_nfc_cfgadvflash_y,
    input              i_nfc_cfgpagesize_y,
    output             o_nfc_cle_a,
    output             o_nfc_nce_a,
    output             o_nfc_nre_a,
    output             o_nfc_nwe_a,
    input              i_nfc_rnb_y,
    input              i_por_reset_y,
    input              i_por_sel_y,
    output             o_sfmc_csn_a,
    input              i_sfmc_sclk_y,
    output             o_sfmc_sclk_a,
    output             o_sfmc_sclk_oe,
    input              i_ssp0_clk_y,
    output             o_ssp0_clk_a,
    output             o_ssp0_clk_oe,
    input              i_ssp0_csn_y,
    output             o_ssp0_csn_a,
    output             o_ssp0_csn_oe,
    input              i_ssp0_rx_y,
    output             o_ssp0_tx_a,
    input              i_ssp1_clk_y,
    output             o_ssp1_clk_a,
    output             o_ssp1_clk_oe,
    input              i_ssp1_csn_y,
    output             o_ssp1_csn_a,
    output             o_ssp1_csn_oe,
    input              i_ssp1_rx_y,
    output             o_ssp1_tx_a,
    input              i_ssp2_clk_y,
    output             o_ssp2_clk_a,
    output             o_ssp2_clk_oe,
    input              i_ssp2_csn_y,
    output             o_ssp2_csn_a,
    output             o_ssp2_csn_oe,
    input              i_ssp2_rx_y,
    output             o_ssp2_tx_a,
    input              i_test_en_y,
    output             o_tg_dvp_h_a,
    output             o_tg_dvp_v_a,
    output             o_tgclk_a,
    input              i_uart0_rxd_y,
    output             o_uart0_txd_a,
    input              i_uart1_rxd_y,
    output             o_uart1_txd_a,
    input              t_aclk,
    input              t_arstn,
    input              t_bist_jtag_tck,
    input              t_bist_jtag_tdi,
    output             t_bist_jtag_tdo,
    output             t_bist_jtag_tdo_oe,
    input              t_bist_jtag_tms,
    input              t_bist_jtag_trst,
    input              t_clk_dvp4,
    input              t_clk_dvp5,
    input              t_clk_dvp6,
    input              t_clk_dvp7,
    input              t_clk_isp0,
    input              t_clk_isp1,
    input              t_clk_isp2,
    input              t_clk_isp3,
    input              t_clk_isp4,
    input              t_clk_isp5,
    input              t_clk_isp6,
    input              t_clk_isp7,
    output             t_ddr_phy_ctrl_div_out_400_a,
    output             t_ddr_phy_ctrl_div_out_800_a,
    output  [  4:  0]  t_ddr_phy_err_a,
    input              t_ddr_phy_ext_ca_cal_en_y,
    output             t_ddr_phy_ext_clock_a,
    input              t_ddr_phy_ext_cmosrcv_y,
    input              t_ddr_phy_ext_dfdqs_y,
    input              t_ddr_phy_ext_en_y,
    output             t_ddr_phy_ext_flock_a,
    input              t_ddr_phy_ext_gatelvl_en_y,
    output             t_ddr_phy_ext_init_complete_a,
    output  [  8:  0]  t_ddr_phy_ext_lock_value_a,
    output             t_ddr_phy_ext_locked_a,
    input   [  3:  0]  t_ddr_phy_ext_mode_y,
    input   [  7:  0]  t_ddr_phy_ext_offsetc_y,
    input              t_ddr_phy_ext_out_y,
    input              t_ddr_phy_ext_rdlvl_en_y,
    input   [  3:  0]  t_ddr_phy_ext_rdlvl_incr_adj_y,
    output  [  3:  0]  t_ddr_phy_ext_rdlvl_vwmc_a,
    input              t_ddr_phy_ext_rdlvl_wr_en_y,
    input              t_ddr_phy_ext_read_y,
    input   [  3:  0]  t_ddr_phy_ext_ref_y,
    input              t_ddr_phy_ext_write_lvl_en_y,
    output             t_ddr_phy_ext_zq_end_a,
    input   [  2:  0]  t_ddr_phy_ext_zq_force_impn_y,
    input   [  2:  0]  t_ddr_phy_ext_zq_force_impp_y,
    input              t_ddr_phy_ext_zq_force_y,
    input   [  2:  0]  t_ddr_phy_ext_zq_mode_dds_y,
    input              t_ddr_phy_highz_y,
    input              t_ddr_phy_mux_y,
    input              t_ddr_phy_nand_y,
    output  [  4:  0]  t_ddr_phy_oky_a,
    input              t_ddr_phy_phy_y,
    input   [  2:  0]  t_ddr_phy_run_y,
    input              t_ddr_phy_scan_y,
    input   [  4:  0]  t_ddr_phy_start_y,
    input              t_ddr_pll_resetb,
    output  [  4:  0]  t_hsp_pll_afc_code,
    output             t_hsp_pll_feed_out,
    output             t_hsp_pll_fout,
    output             t_hsp_pll_lock,
    input              t_hsp_pll_resetb,
    output             t_hsp_pll_sync_m_clk_out,
    output             t_isp0_dvp_clk,
    output             t_isp0_dvp_h,
    output  [ 15:  0]  t_isp0_dvp_p,
    output             t_isp0_dvp_v,
    input              t_isp0_i2cs_scl,
    input              t_isp0_i_i2cs_sda,
    output             t_isp0_o_i2cs_sda,
    output  [  4:  0]  t_isp0_pll_afc_code,
    output             t_isp0_pll_feed_out,
    output             t_isp0_pll_fout,
    output             t_isp0_pll_lock,
    input              t_isp0_pll_resetb,
    output             t_isp0_pll_sync_m_clk_out,
    input              t_isp1_i2cs_scl,
    input              t_isp1_i_i2cs_sda,
    output             t_isp1_o_i2cs_sda,
    output  [  4:  0]  t_isp1_pll_afc_code,
    output             t_isp1_pll_feed_out,
    output             t_isp1_pll_fout,
    output             t_isp1_pll_lock,
    input              t_isp1_pll_resetb,
    output             t_isp1_pll_sync_m_clk_out,
    output             t_isp4_dvp_clk,
    output             t_isp4_dvp_h,
    output  [ 15:  0]  t_isp4_dvp_p,
    output             t_isp4_dvp_v,
    input              t_main_crm_test_rstn,
    output  [  4:  0]  t_main_pll_afc_code,
    output             t_main_pll_feed_out,
    output             t_main_pll_fout,
    output             t_main_pll_lock,
    input              t_main_pll_resetb,
    output             t_main_pll_sync_m_clk_out,
    input   [  1:  0]  t_mipi_rx0_test_sel,
    input   [  1:  0]  t_mipi_rx1_test_sel,
    input              t_mipi_tx_resetb,
    input              t_mtrstn,
    input              t_occ_bypass_pin,
    input              t_occ_reset_pin,
    input              t_occ_test_mode_pin,
    input              t_pll2551_afcini_sel,
    input              t_pll2551_bypass,
    input              t_pll2551_feed_en,
    input              t_pll2551_fout_mask,
    input              t_pll2551_fsel,
    input   [  1:  0]  t_pll2551_icp,
    input   [  1:  0]  t_pll2551_lock_con_dly,
    input   [  1:  0]  t_pll2551_lock_con_in,
    input   [  1:  0]  t_pll2551_lock_con_out,
    input   [  1:  0]  t_pll2551_lock_con_rev,
    input              t_pll2551_lock_en,
    input   [  9:  0]  t_pll2551_m,
    input   [  5:  0]  t_pll2551_p,
    input              t_pll2551_pbias_ctrl,
    input              t_pll2551_pbias_ctrl_en,
    input   [  2:  0]  t_pll2551_s,
    input   [  4:  0]  t_pll2551_tst_afc,
    input              t_pll2551_tst_en,
    input              t_pll2551_vcoini_en,
    output  [  4:  0]  t_pll2651_afc_code,
    input              t_pll2651_afc_enb,
    input              t_pll2651_afcinit_sel,
    input              t_pll2651_bypass,
    input   [  4:  0]  t_pll2651_extafc,
    output             t_pll2651_fout,
    input              t_pll2651_fout_mask,
    input              t_pll2651_fsel,
    input              t_pll2651_fvco_en,
    output             t_pll2651_fvco_out,
    input   [  1:  0]  t_pll2651_icp,
    input   [ 15:  0]  t_pll2651_k,
    input              t_pll2651_lrd_en,
    input   [  8:  0]  t_pll2651_m,
    input   [  7:  0]  t_pll2651_mfr,
    input   [  5:  0]  t_pll2651_mrr,
    input   [  5:  0]  t_pll2651_p,
    input              t_pll2651_pbias_ctrl,
    input              t_pll2651_pbias_ctrl_en,
    input   [  2:  0]  t_pll2651_s,
    input   [  1:  0]  t_pll2651_sel_pf,
    input              t_pll2651_sscg_en,
    input              t_pll2651_vco_boost,
    input              t_pll_sr_ctrl_clk,
    input              t_pll_sr_ctrl_in,
    input              t_pll_sr_ctrl_rst,
    input              t_rstn_isp0,
    input              t_rstn_isp4,
    input              t_scan_cg_en,
    input              t_scan_clk0,
    input              t_scan_clk1,
    input              t_scan_clk2,
    input              t_scan_clk3,
    input              t_scan_clk4,
    input              t_scan_clk5,
    input              t_scan_clk6,
    input              t_scan_comp_en,
    input              t_scan_in00,
    input              t_scan_in01,
    input              t_scan_in02,
    input              t_scan_in03,
    input              t_scan_in04,
    input              t_scan_in05,
    input              t_scan_in06,
    input              t_scan_in07,
    input              t_scan_in08,
    input              t_scan_in09,
    input              t_scan_in10,
    input              t_scan_in11,
    input              t_scan_in12,
    input              t_scan_in13,
    input              t_scan_in14,
    input              t_scan_in15,
    input              t_scan_in16,
    input              t_scan_in17,
    input              t_scan_in18,
    input              t_scan_in19,
    input              t_scan_in20,
    input              t_scan_in21,
    input              t_scan_in22,
    input              t_scan_in23,
    input              t_scan_in24,
    input              t_scan_in25,
    input              t_scan_in26,
    input              t_scan_in27,
    input              t_scan_in28,
    input              t_scan_in29,
    input              t_scan_in30,
    output             t_scan_out00,
    output             t_scan_out01,
    output             t_scan_out02,
    output             t_scan_out03,
    output             t_scan_out04,
    output             t_scan_out05,
    output             t_scan_out06,
    output             t_scan_out07,
    output             t_scan_out08,
    output             t_scan_out09,
    output             t_scan_out10,
    output             t_scan_out11,
    output             t_scan_out12,
    output             t_scan_out13,
    output             t_scan_out14,
    output             t_scan_out15,
    output             t_scan_out16,
    output             t_scan_out17,
    output             t_scan_out18,
    output             t_scan_out19,
    output             t_scan_out20,
    output             t_scan_out21,
    output             t_scan_out22,
    output             t_scan_out23,
    output             t_scan_out24,
    output             t_scan_out25,
    output             t_scan_out26,
    output             t_scan_out27,
    output             t_scan_out28,
    output             t_scan_out29,
    output             t_scan_out30,
    input              t_scan_se,
    input              t_test_rstn,
    input   [ 33:  0]  t_tg_data,
    output  [  4:  0]  t_tg_pll_afc_code,
    output             t_tg_pll_feed_out,
    output             t_tg_pll_fout,
    output             t_tg_pll_lock,
    input              t_tg_pll_resetb,
    output             t_tg_pll_sync_m_clk_out,
    input              t_tgclk,
    input   [  3:  0]  MIPI_DN_RX5,
    inout   [ 31:  0]  DDR_MEM_DQ,
    input   [  3:  0]  MIPI_DP_RX4,
    inout   [  3:  0]  DDR_MEM_DM,
    input   [  3:  0]  MIPI_DN_RX0,
    inout   [  1:  0]  DDR_MEM_CKE,
    inout   [  3:  0]  DDR_MEM_DQS_N,
    input   [  3:  0]  MIPI_DN_RX4,
    input   [  3:  0]  MIPI_DP_RX2,
    inout   [ 15:  0]  DDR_MEM_A,
    inout   [  2:  0]  DDR_MEM_BA,
    output  [  3:  0]  MIPI_DN_TX,
    inout   [  1:  0]  DDR_MEM_ODT,
    output  [  3:  0]  MIPI_DP_TX,
    input   [  3:  0]  MIPI_DP_RX5,
    input   [  3:  0]  MIPI_DP_RX6,
    input   [  3:  0]  MIPI_DN_RX7,
    input   [  3:  0]  MIPI_DP_RX3,
    input   [  3:  0]  MIPI_DP_RX0,
    output  [  3:  0]  MIPI_HS_DO_TX,
    input   [  3:  0]  MIPI_DN_RX3,
    output  [  3:  0]  MIPI_HS_DO_RX0,
    input   [  3:  0]  MIPI_DN_RX2,
    input   [  3:  0]  MIPI_DP_RX1,
    inout   [  1:  0]  DDR_MEM_CSN,
    inout   [  3:  0]  DDR_MEM_DQS_P,
    output  [  3:  0]  MIPI_HS_DO_RX4,
    input   [  3:  0]  MIPI_DN_RX1,
    input   [  3:  0]  MIPI_DP_RX7,
    input   [  3:  0]  MIPI_DN_RX6,
    inout              DDR_MEM_CASN,
    input              DDR_MEM_CKEIN,
    output             DDR_MEM_CK_N,
    output             DDR_MEM_CK_P,
    inout              DDR_MEM_RASN,
    inout              DDR_MEM_RESET_N,
    inout              DDR_MEM_WEN,
    inout              DDR_VREF0,
    inout              DDR_VREF1,
    inout              DDR_ZQ,
    input              MIPI_CHIP_EN_MR0,
    input              MIPI_CHIP_EN_MR1,
    input              MIPI_CHIP_EN_TX,
    input              MIPI_CLKN_RX0,
    input              MIPI_CLKN_RX1,
    input              MIPI_CLKN_RX2,
    input              MIPI_CLKN_RX3,
    input              MIPI_CLKN_RX4,
    input              MIPI_CLKN_RX5,
    input              MIPI_CLKN_RX6,
    input              MIPI_CLKN_RX7,
    output             MIPI_CLKN_TX,
    input              MIPI_CLKP_RX0,
    input              MIPI_CLKP_RX1,
    input              MIPI_CLKP_RX2,
    input              MIPI_CLKP_RX3,
    input              MIPI_CLKP_RX4,
    input              MIPI_CLKP_RX5,
    input              MIPI_CLKP_RX6,
    input              MIPI_CLKP_RX7,
    output             MIPI_CLKP_TX,
    output             MIPI_HS_CKO_RX0,
    output             MIPI_HS_CKO_RX4,
    output             MIPI_HS_CKO_TX,
    output             MIPI_TEST_CLK_A0,
    output             MIPI_TEST_VMON_OUT_RX0,
    output             MIPI_TEST_VMON_OUT_RX4,
    output             MIPI_TEST_VMON_OUT_TX,
    input              i_xin_CK,
    output  [262:  0]  o_core_ds0,
    output  [262:  0]  o_core_ds1,
    output  [262:  0]  o_core_pe,
    output  [262:  0]  o_core_ps,
    output  [262:  0]  o_core_is,
    output  [262:  0]  o_core_sr,
    output  [263:263]  o_core_e0,
    output  [263:263]  o_core_e1,
    output  [263:263]  o_core_sf0,
    output  [263:263]  o_core_sf1,
    output  [262:  0]  o_core_enb,
    input              i_TM_ALL,
    input              i_TM_0_DC,
    input              i_TM_1_NAND,
    input              i_TM_2_SCAN,
    input              i_TM_3_BIST,
    input              i_TM_4_PLL,
    input              i_TM_5_DDR_PHY,
    input              i_TM_6_OCC,
    input              i_TM_7_MIPI_TEST,
    output  [525:  0]  o_func_sel
);




endmodule