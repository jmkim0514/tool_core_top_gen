module peri_hpdf (
    input           i_aclk    ,
    input           i_aresetn ,
    input  [3:0]    i_peri_awid    ,
    input  [31:0]   i_peri_awaddr  ,
    input  [3:0]    i_peri_awlen   ,
    input  [2:0]    i_peri_awsize  ,
    input  [1:0]    i_peri_awburst ,
    input  [1:0]    i_peri_awlock  ,
    input  [3:0]    i_peri_awcache ,
    input  [2:0]    i_peri_awprot  ,
    input           i_peri_awvalid ,
    output          o_peri_awready ,
    input  [3:0]    i_peri_wid     ,
    input  [127:0]  i_peri_wdata   ,
    input  [15:0]   i_peri_wstrb   ,
    input           i_peri_wlast   ,
    input           i_peri_wvalid  ,
    output          o_peri_wready  ,
    output [3:0]    o_peri_bid     ,
    output [1:0]    o_peri_bresp   ,
    output          o_peri_bvalid  ,
    input           i_peri_bready  ,
    input  [3:0]    i_peri_arid    ,
    input  [31:0]   i_peri_araddr  ,
    input  [3:0]    i_peri_arlen   ,
    input  [2:0]    i_peri_arsize  ,
    input  [1:0]    i_peri_arburst ,
    input  [1:0]    i_peri_arlock  ,
    input  [3:0]    i_peri_arcache ,
    input  [2:0]    i_peri_arprot  ,
    input           i_peri_arvalid ,
    output          o_peri_arready ,
    output [3:0]    o_peri_rid     ,
    output [127:0]  o_peri_rdata   ,
    output [1:0]    o_peri_rresp   ,
    output          o_peri_rlast   ,
    output          o_peri_rvalid  ,
    input           i_peri_rready  ,
    input           i_pclk         ,
    input           i_presetn      ,
    output          o_irq          ,
    output          o_psel         ,
    output          o_penable      ,
    output [31:0]   o_paddr        ,
    output          o_pwrite       ,
    output [31:0]   o_pwdata       ,
    output [2:0]    o_pprot        ,
    output [3:0]    o_pstrb        ,
    input  [31:0]   i_prdata       ,
    input           i_pready       ,
    input           i_pslverr      ,
    output          o_irq_wdt       ,
    output          o_irq_pmu       ,
    output          o_irq_otp       
);


endmodule