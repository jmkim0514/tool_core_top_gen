//==============================================================================
//
// Project : PNAI70X
//
// Verilog RTL(Behavioral) model
//
// This confidential and proprietary source code may be used only as authorized
// by a licensing agreement from ALPHAHOLDINGS Limited. The entire notice above
// must be reproduced on all authorized copies and copies may only be made to
// the extent permitted by a licensing agreement from ALPHAHOLDINGS Limited.
//
// COPYRIGHT (C) ALPHAHOLDINGS, inc. 2022
//
//==============================================================================
// File name : peri_hpdf
// Version : v1.0
// Description :
// Simulator : NC Verilog
// Created by : SoC Designer
// Date : 2022-04-19  20:21
//==============================================================================

module peri_hpdf (
    input              i_test_mode,
    input              i_i2s0_bck_y,
    output             o_i2s0_bck_a,
    output             o_i2s0_bck_oe,
    input              i_i2s0_lrck_y,
    output             o_i2s0_lrck_a,
    output             o_i2s0_lrck_oe,
    output             o_i2s0_codck_a,
    output             o_i2s0_codck_oe,
    output             o_i2s0_txdreq,
    input              i_i2s0_txdack,
    output             o_i2s0_rxdreq,
    input              i_i2s0_rxdack,
    input              i_i2s0_rx_y,
    output             o_i2s0_tx_a,
    input              i_i2s1_bck_y,
    output             o_i2s1_bck_a,
    output             o_i2s1_bck_oe,
    input              i_i2s1_lrck_y,
    output             o_i2s1_lrck_a,
    output             o_i2s1_lrck_oe,
    output             o_i2s1_codck_a,
    output             o_i2s1_codck_oe,
    output             o_i2s1_txdreq,
    input              i_i2s1_txdack,
    output             o_i2s1_rxdreq,
    input              i_i2s1_rxdack,
    input              i_i2s1_rx_y,
    output             o_i2s1_tx_a,
    input              i_i2c0_scl_y,
    output             o_i2c0_scl_a,
    output             o_i2c0_scl_oe,
    input              i_i2c0_sda_y,
    output             o_i2c0_sda_a,
    output             o_i2c0_sda_oe,
    output             o_i2c0_int,
    input              i_i2c1_scl_y,
    output             o_i2c1_scl_a,
    output             o_i2c1_scl_oe,
    input              i_i2c1_sda_y,
    output             o_i2c1_sda_a,
    output             o_i2c1_sda_oe,
    output             o_i2c1_int,
    input              i_i2c2_scl_y,
    output             o_i2c2_scl_a,
    output             o_i2c2_scl_oe,
    input              i_i2c2_sda_y,
    output             o_i2c2_sda_a,
    output             o_i2c2_sda_oe,
    output             o_i2c2_int,
    input              i_i2c3_scl_y,
    output             o_i2c3_scl_a,
    output             o_i2c3_scl_oe,
    input              i_i2c3_sda_y,
    output             o_i2c3_sda_a,
    output             o_i2c3_sda_oe,
    output             o_i2c3_int,
    output             o_uart0_txdmasreq,
    output             o_uart0_rxdmasreq,
    output             o_uart0_txdmabreq,
    output             o_uart0_rxdmabreq,
    input              i_uart0_txdmaclr,
    input              i_uart0_rxdmaclr,
    output             o_uart0_intr,
    input              i_uart0_rxd_y,
    output             o_uart0_txd_a,
    output             o_uart1_txdmasreq,
    output             o_uart1_rxdmasreq,
    output             o_uart1_txdmabreq,
    output             o_uart1_rxdmabreq,
    input              i_uart1_txdmaclr,
    input              i_uart1_rxdmaclr,
    output             o_uart1_intr,
    input              i_uart1_rxd_y,
    output             o_uart1_txd_a,
    output             o_uart2_txdmasreq,
    output             o_uart2_rxdmasreq,
    output             o_uart2_txdmabreq,
    output             o_uart2_rxdmabreq,
    input              i_uart2_txdmaclr,
    input              i_uart2_rxdmaclr,
    output             o_uart2_intr,
    input              i_uart2_rxd_y,
    output             o_uart2_txd_a,
    output             o_uart3_txdmasreq,
    output             o_uart3_rxdmasreq,
    output             o_uart3_txdmabreq,
    output             o_uart3_rxdmabreq,
    input              i_uart3_txdmaclr,
    input              i_uart3_rxdmaclr,
    output             o_uart3_intr,
    input              i_uart3_rxd_y,
    output             o_uart3_txd_a,
    output             o_ssp0_intr,
    output             o_ssp0_txdamsreq,
    output             o_ssp0_rxdmasreq,
    output             o_ssp0_txdmabreq,
    output             o_ssp0_rxdmabreq,
    input              i_ssp0_txdmaclr,
    input              i_ssp0_rxdmaclr,
    input              i_ssp0_clk_y,
    output             o_ssp0_clk_a,
    output             o_ssp0_clk_oe,
    input              i_ssp0_csn_y,
    output             o_ssp0_csn_a,
    output             o_ssp0_csn_oe,
    input              i_ssp0_rx_y,
    output             o_ssp0_tx_a,
    output             o_ssp1_intr,
    output             o_ssp1_txdamsreq,
    output             o_ssp1_rxdmasreq,
    output             o_ssp1_txdmabreq,
    output             o_ssp1_rxdmabreq,
    input              i_ssp1_txdmaclr,
    input              i_ssp1_rxdmaclr,
    input              i_ssp1_clk_y,
    output             o_ssp1_clk_a,
    output             o_ssp1_clk_oe,
    input              i_ssp1_csn_y,
    output             o_ssp1_csn_a,
    output             o_ssp1_csn_oe,
    input              i_ssp1_rx_y,
    output             o_ssp1_tx_a,
    output             o_ssp2_intr,
    output             o_ssp2_txdamsreq,
    output             o_ssp2_rxdmasreq,
    output             o_ssp2_txdmabreq,
    output             o_ssp2_rxdmabreq,
    input              i_ssp2_txdmaclr,
    input              i_ssp2_rxdmaclr,
    input              i_ssp2_clk_y,
    output             o_ssp2_clk_a,
    output             o_ssp2_clk_oe,
    input              i_ssp2_csn_y,
    output             o_ssp2_csn_a,
    output             o_ssp2_csn_oe,
    input              i_ssp2_rx_y,
    output             o_ssp2_tx_a,
    output             o_ssp3_intr,
    output             o_ssp3_txdamsreq,
    output             o_ssp3_rxdmasreq,
    output             o_ssp3_txdmabreq,
    output             o_ssp3_rxdmabreq,
    input              i_ssp3_txdmaclr,
    input              i_ssp3_rxdmaclr,
    input              i_ssp3_clk_y,
    output             o_ssp3_clk_a,
    output             o_ssp3_clk_oe,
    input              i_ssp3_csn_y,
    output             o_ssp3_csn_a,
    output             o_ssp3_csn_oe,
    input              i_ssp3_rx_y,
    output             o_ssp3_tx_a,
    output  [  4:  0]  o_timer0_intr,
    output  [  4:  0]  o_timer1_intr,
    output  [  4:  0]  o_timer2_intr,
    output  [  4:  0]  o_timer3_intr,
    output             o_gpio0_intr,
    input   [  7:  0]  i_gpio0_y,
    output  [  7:  0]  o_gpio0_a,
    output  [  7:  0]  o_gpio0_oe,
    output             o_gpio1_intr,
    input   [  7:  0]  i_gpio1_y,
    output  [  7:  0]  o_gpio1_a,
    output  [  7:  0]  o_gpio1_oe,
    output             o_gpio2_intr,
    input   [  7:  0]  i_gpio2_y,
    output  [  7:  0]  o_gpio2_a,
    output  [  7:  0]  o_gpio2_oe,
    output             o_gpio3_intr,
    input   [  7:  0]  i_gpio3_y,
    output  [  7:  0]  o_gpio3_a,
    output  [  7:  0]  o_gpio3_oe,
    output             o_gpio4_intr,
    input   [  7:  0]  i_gpio4_y,
    output  [  7:  0]  o_gpio4_a,
    output  [  7:  0]  o_gpio4_oe,
    output             o_gpio5_intr,
    input   [  7:  0]  i_gpio5_y,
    output  [  7:  0]  o_gpio5_a,
    output  [  7:  0]  o_gpio5_oe,
    output             o_gpio6_intr,
    input   [  7:  0]  i_gpio6_y,
    output  [  7:  0]  o_gpio6_a,
    output  [  7:  0]  o_gpio6_oe,
    output             o_gpio7_intr,
    input   [  7:  0]  i_gpio7_y,
    output  [  7:  0]  o_gpio7_a,
    output  [  7:  0]  o_gpio7_oe,
    output             o_gpio8_intr,
    input   [  7:  0]  i_gpio8_y,
    output  [  7:  0]  o_gpio8_a,
    output  [  7:  0]  o_gpio8_oe,
    output             o_gpio9_intr,
    input   [  7:  0]  i_gpio9_y,
    output  [  7:  0]  o_gpio9_a,
    output  [  7:  0]  o_gpio9_oe,
    output             o_gpio10_intr,
    input   [  7:  0]  i_gpio10_y,
    output  [  7:  0]  o_gpio10_a,
    output  [  7:  0]  o_gpio10_oe,
    output             o_gpio11_intr,
    input   [  7:  0]  i_gpio11_y,
    output  [  7:  0]  o_gpio11_a,
    output  [  7:  0]  o_gpio11_oe,
    output             o_gpio12_intr,
    input   [  7:  0]  i_gpio12_y,
    output  [  7:  0]  o_gpio12_a,
    output  [  7:  0]  o_gpio12_oe,
    output             o_gpio13_intr,
    input   [  7:  0]  i_gpio13_y,
    output  [  7:  0]  o_gpio13_a,
    output  [  7:  0]  o_gpio13_oe,
    output             o_gpio14_intr,
    input   [  7:  0]  i_gpio14_y,
    output  [  7:  0]  o_gpio14_a,
    output  [  7:  0]  o_gpio14_oe,
    output             o_gpio15_intr,
    input   [  7:  0]  i_gpio15_y,
    output  [  7:  0]  o_gpio15_a,
    output  [  7:  0]  o_gpio15_oe,
    output             o_gpio16_intr,
    input   [  7:  0]  i_gpio16_y,
    output  [  7:  0]  o_gpio16_a,
    output  [  7:  0]  o_gpio16_oe,
    output             o_gpio17_intr,
    input   [  7:  0]  i_gpio17_y,
    output  [  7:  0]  o_gpio17_a,
    output  [  7:  0]  o_gpio17_oe,
    output             o_gpio18_intr,
    input   [  7:  0]  i_gpio18_y,
    output  [  7:  0]  o_gpio18_a,
    output  [  7:  0]  o_gpio18_oe,
    output             o_gpio19_intr,
    input   [  7:  0]  i_gpio19_y,
    output  [  7:  0]  o_gpio19_a,
    output  [  7:  0]  o_gpio19_oe,
    output             o_wdt_intr,
    output             o_wdt_nresetout,
    output             o_rtc_tic_irq0,
    output             o_rtc_tic_irq1,
    output             o_rtc_alarm_irq,
    input              i_rtc_xin_ck,
    output             o_adc_clk,
    output             o_adc_pd,
    output             o_adc_soc,
    output  [  3:  0]  o_adc_sel,
    input              i_adc_eoc,
    input   [ 11:  0]  i_adc_data,
    input              i_clk_peri_hpdf,
    input              i_rstn_peri_hpdf,
    input              i_clk_peri_codec,
    input              i_i2s0_codck_y,
    input              i_i2s1_codck_y,
    output             i_clk_peri_bus,
    output             i_rstn_peri_bus,
    input              i_test_clk,
    input   [  4:  0]  i_cpu_awid_m4_cpu2_peri,
    input   [ 31:  0]  i_cpu_awaddr_m4_cpu2_peri,
    input   [  7:  0]  i_cpu_awlen_m4_cpu2_peri,
    input   [  2:  0]  i_cpu_awsize_m4_cpu2_peri,
    input   [  1:  0]  i_cpu_awburst_m4_cpu2_peri,
    input              i_cpu_awlock_m4_cpu2_peri,
    input   [  3:  0]  i_cpu_awcache_m4_cpu2_peri,
    input   [  2:  0]  i_cpu_awprot_m4_cpu2_peri,
    input              i_cpu_awvalid_m4_cpu2_peri,
    output             o_cpu_awready_m4_cpu2_peri,
    input   [  4:  0]  i_cpu_arid_m4_cpu2_peri,
    input   [ 31:  0]  i_cpu_araddr_m4_cpu2_peri,
    input   [  7:  0]  i_cpu_arlen_m4_cpu2_peri,
    input   [  2:  0]  i_cpu_arsize_m4_cpu2_peri,
    input   [  1:  0]  i_cpu_arburst_m4_cpu2_peri,
    input              i_cpu_arlock_m4_cpu2_peri,
    input   [  3:  0]  i_cpu_arcache_m4_cpu2_peri,
    input   [  2:  0]  i_cpu_arprot_m4_cpu2_peri,
    input              i_cpu_arvalid_m4_cpu2_peri,
    output             o_cpu_arready_m4_cpu2_peri,
    input   [ 31:  0]  i_cpu_wdata_m4_cpu2_peri,
    input   [  3:  0]  i_cpu_wstrb_m4_cpu2_peri,
    input              i_cpu_wlast_m4_cpu2_peri,
    input              i_cpu_wvalid_m4_cpu2_peri,
    output             o_cpu_wready_m4_cpu2_peri,
    output  [  4:  0]  o_cpu_bid_m4_cpu2_peri,
    output  [  1:  0]  o_cpu_bresp_m4_cpu2_peri,
    output             o_cpu_bvalid_m4_cpu2_peri,
    input              i_cpu_bready_m4_cpu2_peri,
    output  [  4:  0]  o_cpu_rid_m4_cpu2_peri,
    output  [  1:  0]  o_cpu_rresp_m4_cpu2_peri,
    output  [ 31:  0]  o_cpu_rdata_m4_cpu2_peri,
    output             o_cpu_rlast_m4_cpu2_peri,
    output             o_cpu_rvalid_m4_cpu2_peri,
    input              i_cpu_rready_m4_cpu2_peri,
    output             o_peri_pselx_codec_hpdf_m3,
    output             o_peri_penable_codec_hpdf_m3,
    output  [ 31:  0]  o_peri_paddr_codec_hpdf_m3,
    output             o_peri_pwrite_codec_hpdf_m3,
    output  [ 31:  0]  o_peri_pwdata_codec_hpdf_m3,
    input   [ 31:  0]  i_peri_prdata_codec_hpdf_m3,
    input              i_peri_pready_codec_hpdf_m3,
    input              i_peri_pslverr_codec_hpdf_m3,
    output             o_peri_pselx_disp_hpdf_m5,
    output             o_peri_penable_disp_hpdf_m5,
    output  [ 31:  0]  o_peri_paddr_disp_hpdf_m5,
    output             o_peri_pwrite_disp_hpdf_m5,
    output  [ 31:  0]  o_peri_pwdata_disp_hpdf_m5,
    input   [ 31:  0]  i_peri_prdata_disp_hpdf_m5,
    input              i_peri_pready_disp_hpdf_m5,
    input              i_peri_pslverr_disp_hpdf_m5,
    output             o_peri_pselx_hsp_hpdf_m2,
    output             o_peri_penable_hsp_hpdf_m2,
    output  [ 31:  0]  o_peri_paddr_hsp_hpdf_m2,
    output             o_peri_pwrite_hsp_hpdf_m2,
    output  [ 31:  0]  o_peri_pwdata_hsp_hpdf_m2,
    input   [ 31:  0]  i_peri_prdata_hsp_hpdf_m2,
    input              i_peri_pready_hsp_hpdf_m2,
    input              i_peri_pslverr_hsp_hpdf_m2,
    output             o_peri_pselx_npu_hpdf_m4,
    output             o_peri_penable_npu_hpdf_m4,
    output  [ 31:  0]  o_peri_paddr_npu_hpdf_m4,
    output             o_peri_pwrite_npu_hpdf_m4,
    output  [ 31:  0]  o_peri_pwdata_npu_hpdf_m4,
    input   [ 31:  0]  i_peri_prdata_npu_hpdf_m4,
    input              i_peri_pready_npu_hpdf_m4,
    input              i_peri_pslverr_npu_hpdf_m4
);

    wire    [33:0]  NC_in;
    wire    [66:0]  NC_out;
    wire    [31:0]  peri_paddr_peri0_m0;
    wire            peri_pselx_peri0_m0;
    wire            peri_penable_peri0_m0;
    wire            peri_pwrite_peri0_m0;
    wire    [31:0]  peri_prdata_peri0_m0;
    wire    [31:0]  peri_pwdata_peri0_m0;
    wire            peri_pready_peri0_m0;
    wire            peri_pslverr_peri0_m0;
    wire            peri_sub_o_crm_apb_psel;
    wire            peri_sub_o_crm_apb_penable;
    wire            peri_sub_o_crm_apb_pwrite;
    wire    [11:0]  peri_sub_o_crm_apb_paddr;
    wire    [31:0]  peri_sub_o_crm_apb_pwdata;
    wire    [31:0]  peri_sub_i_crm_apb_prdata;
    wire            crm_peri_o_clk_pclk_i2s0;
    wire            crm_peri_o_rstn_pclk_i2s0;
    wire            crm_peri_o_clk_pclk_i2s1;
    wire            crm_peri_o_rstn_pclk_i2s1;
    wire            crm_peri_o_clk_pclk_i2c0;
    wire            crm_peri_o_rstn_pclk_i2c0;
    wire            crm_peri_o_clk_pclk_i2c1;
    wire            crm_peri_o_rstn_pclk_i2c1;
    wire            crm_peri_o_clk_pclk_i2c2;
    wire            crm_peri_o_rstn_pclk_i2c2;
    wire            crm_peri_o_clk_pclk_i2c3;
    wire            crm_peri_o_rstn_pclk_i2c3;
    wire            crm_peri_o_clk_pclk_uart0;
    wire            crm_peri_o_rstn_pclk_uart0;
    wire            crm_peri_o_clk_pclk_uart1;
    wire            crm_peri_o_rstn_pclk_uart1;
    wire            crm_peri_o_clk_pclk_uart2;
    wire            crm_peri_o_rstn_pclk_uart2;
    wire            crm_peri_o_clk_pclk_uart3;
    wire            crm_peri_o_rstn_pclk_uart3;
    wire            crm_peri_o_clk_pclk_spi0;
    wire            crm_peri_o_rstn_pclk_spi0;
    wire            crm_peri_o_clk_pclk_spi1;
    wire            crm_peri_o_rstn_pclk_spi1;
    wire            crm_peri_o_clk_pclk_spi2;
    wire            crm_peri_o_rstn_pclk_spi2;
    wire            crm_peri_o_clk_pclk_spi3;
    wire            crm_peri_o_rstn_pclk_spi3;
    wire            crm_peri_o_clk_pclk_timer0;
    wire            crm_peri_o_rstn_pclk_timer0;
    wire            crm_peri_o_clk_pclk_timer1;
    wire            crm_peri_o_rstn_pclk_timer1;
    wire            crm_peri_o_clk_pclk_timer2;
    wire            crm_peri_o_rstn_pclk_timer2;
    wire            crm_peri_o_clk_pclk_timer3;
    wire            crm_peri_o_rstn_pclk_timer3;
    wire            crm_peri_o_clk_pclk_gpio0;
    wire            crm_peri_o_rstn_pclk_gpio0;
    wire            crm_peri_o_clk_pclk_gpio1;
    wire            crm_peri_o_rstn_pclk_gpio1;
    wire            crm_peri_o_clk_pclk_gpio2;
    wire            crm_peri_o_rstn_pclk_gpio2;
    wire            crm_peri_o_clk_pclk_gpio3;
    wire            crm_peri_o_rstn_pclk_gpio3;
    wire            crm_peri_o_clk_pclk_gpio4;
    wire            crm_peri_o_rstn_pclk_gpio4;
    wire            crm_peri_o_clk_pclk_gpio5;
    wire            crm_peri_o_rstn_pclk_gpio5;
    wire            crm_peri_o_clk_pclk_gpio6;
    wire            crm_peri_o_rstn_pclk_gpio6;
    wire            crm_peri_o_clk_pclk_gpio7;
    wire            crm_peri_o_rstn_pclk_gpio7;
    wire            crm_peri_o_clk_pclk_gpio8;
    wire            crm_peri_o_rstn_pclk_gpio8;
    wire            crm_peri_o_clk_pclk_gpio9;
    wire            crm_peri_o_rstn_pclk_gpio9;
    wire            crm_peri_o_clk_pclk_gpio10;
    wire            crm_peri_o_rstn_pclk_gpio10;
    wire            crm_peri_o_clk_pclk_gpio11;
    wire            crm_peri_o_rstn_pclk_gpio11;
    wire            crm_peri_o_clk_pclk_gpio12;
    wire            crm_peri_o_rstn_pclk_gpio12;
    wire            crm_peri_o_clk_pclk_gpio13;
    wire            crm_peri_o_rstn_pclk_gpio13;
    wire            crm_peri_o_clk_pclk_gpio14;
    wire            crm_peri_o_rstn_pclk_gpio14;
    wire            crm_peri_o_clk_pclk_gpio15;
    wire            crm_peri_o_rstn_pclk_gpio15;
    wire            crm_peri_o_clk_pclk_gpio16;
    wire            crm_peri_o_rstn_pclk_gpio16;
    wire            crm_peri_o_clk_pclk_gpio17;
    wire            crm_peri_o_rstn_pclk_gpio17;
    wire            crm_peri_o_clk_pclk_gpio18;
    wire            crm_peri_o_rstn_pclk_gpio18;
    wire            crm_peri_o_clk_pclk_gpio19;
    wire            crm_peri_o_rstn_pclk_gpio19;
    wire            crm_peri_o_clk_pclk_wdt;
    wire            crm_peri_o_rstn_pclk_wdt;
    wire            crm_peri_o_clk_pclk_rtc;
    wire            crm_peri_o_rstn_pclk_rtc;
    wire            crm_peri_o_clk_pclk_adc;
    wire            crm_peri_o_rstn_pclk_adc;
    wire            crm_peri_o_clk_peri_bus;
    wire            crm_peri_o_rstn_peri_bus;
    wire            crm_peri_o_clk_codec_clk0;
    wire            crm_peri_o_clk_codec_clk1;

    assign  i_clk_peri_bus = crm_peri_o_clk_peri_bus;
    assign  i_rstn_peri_bus = crm_peri_o_rstn_peri_bus;

    nic400_peri_bus_r0p00 u_peri_bus (
        .paddr_codec_hpdf_m3     (o_peri_paddr_codec_hpdf_m3),
        .pselx_codec_hpdf_m3     (o_peri_pselx_codec_hpdf_m3),
        .penable_codec_hpdf_m3   (o_peri_penable_codec_hpdf_m3),
        .pwrite_codec_hpdf_m3    (o_peri_pwrite_codec_hpdf_m3),
        .prdata_codec_hpdf_m3    (i_peri_prdata_codec_hpdf_m3),
        .pwdata_codec_hpdf_m3    (o_peri_pwdata_codec_hpdf_m3),
        .pready_codec_hpdf_m3    (i_peri_pready_codec_hpdf_m3),
        .pslverr_codec_hpdf_m3   (i_peri_pslverr_codec_hpdf_m3),
        .awid_cpu2peri_s0        (i_cpu_awid_m4_cpu2_peri),
        .awaddr_cpu2peri_s0      (i_cpu_awaddr_m4_cpu2_peri),
        .awlen_cpu2peri_s0       (i_cpu_awlen_m4_cpu2_peri),
        .awsize_cpu2peri_s0      (i_cpu_awsize_m4_cpu2_peri),
        .awburst_cpu2peri_s0     (i_cpu_awburst_m4_cpu2_peri),
        .awlock_cpu2peri_s0      (i_cpu_awlock_m4_cpu2_peri),
        .awcache_cpu2peri_s0     (i_cpu_awcache_m4_cpu2_peri),
        .awprot_cpu2peri_s0      (i_cpu_awprot_m4_cpu2_peri),
        .awvalid_cpu2peri_s0     (i_cpu_awvalid_m4_cpu2_peri),
        .awready_cpu2peri_s0     (o_cpu_awready_m4_cpu2_peri),
        .wdata_cpu2peri_s0       (i_cpu_wdata_m4_cpu2_peri),
        .wstrb_cpu2peri_s0       (i_cpu_wstrb_m4_cpu2_peri),
        .wlast_cpu2peri_s0       (i_cpu_wlast_m4_cpu2_peri),
        .wvalid_cpu2peri_s0      (i_cpu_wvalid_m4_cpu2_peri),
        .wready_cpu2peri_s0      (o_cpu_wready_m4_cpu2_peri),
        .bid_cpu2peri_s0         (o_cpu_bid_m4_cpu2_peri),
        .bresp_cpu2peri_s0       (o_cpu_bresp_m4_cpu2_peri),
        .bvalid_cpu2peri_s0      (o_cpu_bvalid_m4_cpu2_peri),
        .bready_cpu2peri_s0      (i_cpu_bready_m4_cpu2_peri),
        .arid_cpu2peri_s0        (i_cpu_arid_m4_cpu2_peri),
        .araddr_cpu2peri_s0      (i_cpu_araddr_m4_cpu2_peri),
        .arlen_cpu2peri_s0       (i_cpu_arlen_m4_cpu2_peri),
        .arsize_cpu2peri_s0      (i_cpu_arsize_m4_cpu2_peri),
        .arburst_cpu2peri_s0     (i_cpu_arburst_m4_cpu2_peri),
        .arlock_cpu2peri_s0      (i_cpu_arlock_m4_cpu2_peri),
        .arcache_cpu2peri_s0     (i_cpu_arcache_m4_cpu2_peri),
        .arprot_cpu2peri_s0      (i_cpu_arprot_m4_cpu2_peri),
        .arvalid_cpu2peri_s0     (i_cpu_arvalid_m4_cpu2_peri),
        .arready_cpu2peri_s0     (o_cpu_arready_m4_cpu2_peri),
        .rid_cpu2peri_s0         (o_cpu_rid_m4_cpu2_peri),
        .rdata_cpu2peri_s0       (o_cpu_rdata_m4_cpu2_peri),
        .rresp_cpu2peri_s0       (o_cpu_rresp_m4_cpu2_peri),
        .rlast_cpu2peri_s0       (o_cpu_rlast_m4_cpu2_peri),
        .rvalid_cpu2peri_s0      (o_cpu_rvalid_m4_cpu2_peri),
        .rready_cpu2peri_s0      (i_cpu_rready_m4_cpu2_peri),
        .paddr_ddr_hpdf_m6       (NC_out[31:0]),
        .pselx_ddr_hpdf_m6       (NC_out[32]),
        .penable_ddr_hpdf_m6     (NC_out[33]),
        .pwrite_ddr_hpdf_m6      (NC_out[34]),
        .prdata_ddr_hpdf_m6      (NC_in[31:0]),
        .pwdata_ddr_hpdf_m6      (NC_out[66:35]),
        .pready_ddr_hpdf_m6      (NC_in[32]),
        .pslverr_ddr_hpdf_m6     (NC_in[33]),
        .paddr_disp_hpdf_m5      (o_peri_paddr_disp_hpdf_m5),
        .pselx_disp_hpdf_m5      (o_peri_pselx_disp_hpdf_m5),
        .penable_disp_hpdf_m5    (o_peri_penable_disp_hpdf_m5),
        .pwrite_disp_hpdf_m5     (o_peri_pwrite_disp_hpdf_m5),
        .prdata_disp_hpdf_m5     (i_peri_prdata_disp_hpdf_m5),
        .pwdata_disp_hpdf_m5     (o_peri_pwdata_disp_hpdf_m5),
        .pready_disp_hpdf_m5     (i_peri_pready_disp_hpdf_m5),
        .pslverr_disp_hpdf_m5    (i_peri_pslverr_disp_hpdf_m5),
        .paddr_hsp_hpdf_m2       (o_peri_paddr_hsp_hpdf_m2),
        .pselx_hsp_hpdf_m2       (o_peri_pselx_hsp_hpdf_m2),
        .penable_hsp_hpdf_m2     (o_peri_penable_hsp_hpdf_m2),
        .pwrite_hsp_hpdf_m2      (o_peri_pwrite_hsp_hpdf_m2),
        .prdata_hsp_hpdf_m2      (i_peri_prdata_hsp_hpdf_m2),
        .pwdata_hsp_hpdf_m2      (o_peri_pwdata_hsp_hpdf_m2),
        .pready_hsp_hpdf_m2      (i_peri_pready_hsp_hpdf_m2),
        .pslverr_hsp_hpdf_m2     (i_peri_pslverr_hsp_hpdf_m2),
        .paddr_npu_hpdf_m4       (o_peri_paddr_npu_hpdf_m4),
        .pselx_npu_hpdf_m4       (o_peri_pselx_npu_hpdf_m4),
        .penable_npu_hpdf_m4     (o_peri_penable_npu_hpdf_m4),
        .pwrite_npu_hpdf_m4      (o_peri_pwrite_npu_hpdf_m4),
        .prdata_npu_hpdf_m4      (i_peri_prdata_npu_hpdf_m4),
        .pwdata_npu_hpdf_m4      (o_peri_pwdata_npu_hpdf_m4),
        .pready_npu_hpdf_m4      (i_peri_pready_npu_hpdf_m4),
        .pslverr_npu_hpdf_m4     (i_peri_pslverr_npu_hpdf_m4),
        .paddr_peri0_m0          (peri_paddr_peri0_m0),
        .pselx_peri0_m0          (peri_pselx_peri0_m0),
        .penable_peri0_m0        (peri_penable_peri0_m0),
        .pwrite_peri0_m0         (peri_pwrite_peri0_m0),
        .prdata_peri0_m0         (peri_prdata_peri0_m0),
        .pwdata_peri0_m0         (peri_pwdata_peri0_m0),
        .pready_peri0_m0         (peri_pready_peri0_m0),
        .pslverr_peri0_m0        (peri_pslverr_peri0_m0),
        .mainclk                 (crm_peri_o_clk_peri_bus),
        .mainclk_r               (crm_peri_o_clk_peri_bus),
        .mainclken               (1'h1),
        .mainresetn              (crm_peri_o_rstn_peri_bus),
        .mainresetn_r            (crm_peri_o_rstn_peri_bus)
    );

    peri_sub u_peri_sub (
        .i_paddr_peri0_m0        (peri_paddr_peri0_m0),
        .i_pselx_peri0_m0        (peri_pselx_peri0_m0),
        .i_penable_peri0_m0      (peri_penable_peri0_m0),
        .i_pwrite_peri0_m0       (peri_pwrite_peri0_m0),
        .o_prdata_peri0_m0       (peri_prdata_peri0_m0),
        .i_pwdata_peri0_m0       (peri_pwdata_peri0_m0),
        .o_pready_peri0_m0       (peri_pready_peri0_m0),
        .o_pslverr_peri0_m0      (peri_pslverr_peri0_m0),
        .o_crm_apb_psel          (peri_sub_o_crm_apb_psel),
        .o_crm_apb_penable       (peri_sub_o_crm_apb_penable),
        .o_crm_apb_pwrite        (peri_sub_o_crm_apb_pwrite),
        .o_crm_apb_paddr         (peri_sub_o_crm_apb_paddr),
        .o_crm_apb_pwdata        (peri_sub_o_crm_apb_pwdata),
        .i_crm_apb_prdata        (peri_sub_i_crm_apb_prdata),
        .i_clk_pclk_i2s0         (crm_peri_o_clk_pclk_i2s0),
        .i_rstn_pclk_i2s0        (crm_peri_o_rstn_pclk_i2s0),
        .i_clk_pclk_i2s1         (crm_peri_o_clk_pclk_i2s1),
        .i_rstn_pclk_i2s1        (crm_peri_o_rstn_pclk_i2s1),
        .i_clk_pclk_i2c0         (crm_peri_o_clk_pclk_i2c0),
        .i_rstn_pclk_i2c0        (crm_peri_o_rstn_pclk_i2c0),
        .i_clk_pclk_i2c1         (crm_peri_o_clk_pclk_i2c1),
        .i_rstn_pclk_i2c1        (crm_peri_o_rstn_pclk_i2c1),
        .i_clk_pclk_i2c2         (crm_peri_o_clk_pclk_i2c2),
        .i_rstn_pclk_i2c2        (crm_peri_o_rstn_pclk_i2c2),
        .i_clk_pclk_i2c3         (crm_peri_o_clk_pclk_i2c3),
        .i_rstn_pclk_i2c3        (crm_peri_o_rstn_pclk_i2c3),
        .i_clk_pclk_uart0        (crm_peri_o_clk_pclk_uart0),
        .i_rstn_pclk_uart0       (crm_peri_o_rstn_pclk_uart0),
        .i_clk_pclk_uart1        (crm_peri_o_clk_pclk_uart1),
        .i_rstn_pclk_uart1       (crm_peri_o_rstn_pclk_uart1),
        .i_clk_pclk_uart2        (crm_peri_o_clk_pclk_uart2),
        .i_rstn_pclk_uart2       (crm_peri_o_rstn_pclk_uart2),
        .i_clk_pclk_uart3        (crm_peri_o_clk_pclk_uart3),
        .i_rstn_pclk_uart3       (crm_peri_o_rstn_pclk_uart3),
        .i_clk_pclk_spi0         (crm_peri_o_clk_pclk_spi0),
        .i_rstn_pclk_spi0        (crm_peri_o_rstn_pclk_spi0),
        .i_clk_pclk_spi1         (crm_peri_o_clk_pclk_spi1),
        .i_rstn_pclk_spi1        (crm_peri_o_rstn_pclk_spi1),
        .i_clk_pclk_spi2         (crm_peri_o_clk_pclk_spi2),
        .i_rstn_pclk_spi2        (crm_peri_o_rstn_pclk_spi2),
        .i_clk_pclk_spi3         (crm_peri_o_clk_pclk_spi3),
        .i_rstn_pclk_spi3        (crm_peri_o_rstn_pclk_spi3),
        .i_clk_pclk_timer0       (crm_peri_o_clk_pclk_timer0),
        .i_rstn_pclk_timer0      (crm_peri_o_rstn_pclk_timer0),
        .i_clk_pclk_timer1       (crm_peri_o_clk_pclk_timer1),
        .i_rstn_pclk_timer1      (crm_peri_o_rstn_pclk_timer1),
        .i_clk_pclk_timer2       (crm_peri_o_clk_pclk_timer2),
        .i_rstn_pclk_timer2      (crm_peri_o_rstn_pclk_timer2),
        .i_clk_pclk_timer3       (crm_peri_o_clk_pclk_timer3),
        .i_rstn_pclk_timer3      (crm_peri_o_rstn_pclk_timer3),
        .i_clk_pclk_gpio0        (crm_peri_o_clk_pclk_gpio0),
        .i_rstn_pclk_gpio0       (crm_peri_o_rstn_pclk_gpio0),
        .i_clk_pclk_gpio1        (crm_peri_o_clk_pclk_gpio1),
        .i_rstn_pclk_gpio1       (crm_peri_o_rstn_pclk_gpio1),
        .i_clk_pclk_gpio2        (crm_peri_o_clk_pclk_gpio2),
        .i_rstn_pclk_gpio2       (crm_peri_o_rstn_pclk_gpio2),
        .i_clk_pclk_gpio3        (crm_peri_o_clk_pclk_gpio3),
        .i_rstn_pclk_gpio3       (crm_peri_o_rstn_pclk_gpio3),
        .i_clk_pclk_gpio4        (crm_peri_o_clk_pclk_gpio4),
        .i_rstn_pclk_gpio4       (crm_peri_o_rstn_pclk_gpio4),
        .i_clk_pclk_gpio5        (crm_peri_o_clk_pclk_gpio5),
        .i_rstn_pclk_gpio5       (crm_peri_o_rstn_pclk_gpio5),
        .i_clk_pclk_gpio6        (crm_peri_o_clk_pclk_gpio6),
        .i_rstn_pclk_gpio6       (crm_peri_o_rstn_pclk_gpio6),
        .i_clk_pclk_gpio7        (crm_peri_o_clk_pclk_gpio7),
        .i_rstn_pclk_gpio7       (crm_peri_o_rstn_pclk_gpio7),
        .i_clk_pclk_gpio8        (crm_peri_o_clk_pclk_gpio8),
        .i_rstn_pclk_gpio8       (crm_peri_o_rstn_pclk_gpio8),
        .i_clk_pclk_gpio9        (crm_peri_o_clk_pclk_gpio9),
        .i_rstn_pclk_gpio9       (crm_peri_o_rstn_pclk_gpio9),
        .i_clk_pclk_gpio10       (crm_peri_o_clk_pclk_gpio10),
        .i_rstn_pclk_gpio10      (crm_peri_o_rstn_pclk_gpio10),
        .i_clk_pclk_gpio11       (crm_peri_o_clk_pclk_gpio11),
        .i_rstn_pclk_gpio11      (crm_peri_o_rstn_pclk_gpio11),
        .i_clk_pclk_gpio12       (crm_peri_o_clk_pclk_gpio12),
        .i_rstn_pclk_gpio12      (crm_peri_o_rstn_pclk_gpio12),
        .i_clk_pclk_gpio13       (crm_peri_o_clk_pclk_gpio13),
        .i_rstn_pclk_gpio13      (crm_peri_o_rstn_pclk_gpio13),
        .i_clk_pclk_gpio14       (crm_peri_o_clk_pclk_gpio14),
        .i_rstn_pclk_gpio14      (crm_peri_o_rstn_pclk_gpio14),
        .i_clk_pclk_gpio15       (crm_peri_o_clk_pclk_gpio15),
        .i_rstn_pclk_gpio15      (crm_peri_o_rstn_pclk_gpio15),
        .i_clk_pclk_gpio16       (crm_peri_o_clk_pclk_gpio16),
        .i_rstn_pclk_gpio16      (crm_peri_o_rstn_pclk_gpio16),
        .i_clk_pclk_gpio17       (crm_peri_o_clk_pclk_gpio17),
        .i_rstn_pclk_gpio17      (crm_peri_o_rstn_pclk_gpio17),
        .i_clk_pclk_gpio18       (crm_peri_o_clk_pclk_gpio18),
        .i_rstn_pclk_gpio18      (crm_peri_o_rstn_pclk_gpio18),
        .i_clk_pclk_gpio19       (crm_peri_o_clk_pclk_gpio19),
        .i_rstn_pclk_gpio19      (crm_peri_o_rstn_pclk_gpio19),
        .i_clk_pclk_wdt          (crm_peri_o_clk_pclk_wdt),
        .i_rstn_pclk_wdt         (crm_peri_o_rstn_pclk_wdt),
        .i_clk_pclk_rtc          (crm_peri_o_clk_pclk_rtc),
        .i_rstn_pclk_rtc         (crm_peri_o_rstn_pclk_rtc),
        .i_clk_pclk_adc          (crm_peri_o_clk_pclk_adc),
        .i_rstn_pclk_adc         (crm_peri_o_rstn_pclk_adc),
        .i_clk_peri_bus          (crm_peri_o_clk_peri_bus),
        .i_rstn_peri_bus         (crm_peri_o_rstn_peri_bus),
        .i_scan_tmode            (i_test_mode),
        .i_i2s0_bck_y            (i_i2s0_bck_y),
        .o_i2s0_bck_a            (o_i2s0_bck_a),
        .o_i2s0_bck_oe           (o_i2s0_bck_oe),
        .i_i2s0_lrck_y           (i_i2s0_lrck_y),
        .o_i2s0_lrck_a           (o_i2s0_lrck_a),
        .o_i2s0_lrck_oe          (o_i2s0_lrck_oe),
        .i_i2s0_codck_y          (crm_peri_o_clk_codec_clk0),
        .o_i2s0_codck_a          (o_i2s0_codck_a),
        .o_i2s0_codck_oe         (o_i2s0_codck_oe),
        .o_i2s0_txdreq           (o_i2s0_txdreq),
        .i_i2s0_txdack           (i_i2s0_txdack),
        .o_i2s0_rxdreq           (o_i2s0_rxdreq),
        .i_i2s0_rxdack           (i_i2s0_rxdack),
        .i_i2s0_rx_y             (i_i2s0_rx_y),
        .o_i2s0_tx_a             (o_i2s0_tx_a),
        .i_i2s1_bck_y            (i_i2s1_bck_y),
        .o_i2s1_bck_a            (o_i2s1_bck_a),
        .o_i2s1_bck_oe           (o_i2s1_bck_oe),
        .i_i2s1_lrck_y           (i_i2s1_lrck_y),
        .o_i2s1_lrck_a           (o_i2s1_lrck_a),
        .o_i2s1_lrck_oe          (o_i2s1_lrck_oe),
        .i_i2s1_codck_y          (crm_peri_o_clk_codec_clk1),
        .o_i2s1_codck_a          (o_i2s1_codck_a),
        .o_i2s1_codck_oe         (o_i2s1_codck_oe),
        .o_i2s1_txdreq           (o_i2s1_txdreq),
        .i_i2s1_txdack           (i_i2s1_txdack),
        .o_i2s1_rxdreq           (o_i2s1_rxdreq),
        .i_i2s1_rxdack           (i_i2s1_rxdack),
        .i_i2s1_rx_y             (i_i2s1_rx_y),
        .o_i2s1_tx_a             (o_i2s1_tx_a),
        .i_i2c0_scl_y            (i_i2c0_scl_y),
        .o_i2c0_scl_a            (o_i2c0_scl_a),
        .o_i2c0_scl_oe           (o_i2c0_scl_oe),
        .i_i2c0_sda_y            (i_i2c0_sda_y),
        .o_i2c0_sda_a            (o_i2c0_sda_a),
        .o_i2c0_sda_oe           (o_i2c0_sda_oe),
        .o_i2c0_int              (o_i2c0_int),
        .i_i2c1_scl_y            (i_i2c1_scl_y),
        .o_i2c1_scl_a            (o_i2c1_scl_a),
        .o_i2c1_scl_oe           (o_i2c1_scl_oe),
        .i_i2c1_sda_y            (i_i2c1_sda_y),
        .o_i2c1_sda_a            (o_i2c1_sda_a),
        .o_i2c1_sda_oe           (o_i2c1_sda_oe),
        .o_i2c1_int              (o_i2c1_int),
        .i_i2c2_scl_y            (i_i2c2_scl_y),
        .o_i2c2_scl_a            (o_i2c2_scl_a),
        .o_i2c2_scl_oe           (o_i2c2_scl_oe),
        .i_i2c2_sda_y            (i_i2c2_sda_y),
        .o_i2c2_sda_a            (o_i2c2_sda_a),
        .o_i2c2_sda_oe           (o_i2c2_sda_oe),
        .o_i2c2_int              (o_i2c2_int),
        .i_i2c3_scl_y            (i_i2c3_scl_y),
        .o_i2c3_scl_a            (o_i2c3_scl_a),
        .o_i2c3_scl_oe           (o_i2c3_scl_oe),
        .i_i2c3_sda_y            (i_i2c3_sda_y),
        .o_i2c3_sda_a            (o_i2c3_sda_a),
        .o_i2c3_sda_oe           (o_i2c3_sda_oe),
        .o_i2c3_int              (o_i2c3_int),
        .o_uart0_txdmasreq       (o_uart0_txdmasreq),
        .o_uart0_rxdmasreq       (o_uart0_rxdmasreq),
        .o_uart0_txdmabreq       (o_uart0_txdmabreq),
        .o_uart0_rxdmabreq       (o_uart0_rxdmabreq),
        .i_uart0_txdmaclr        (i_uart0_txdmaclr),
        .i_uart0_rxdmaclr        (i_uart0_rxdmaclr),
        .o_uart0_intr            (o_uart0_intr),
        .i_uart0_rxd_y           (i_uart0_rxd_y),
        .o_uart0_txd_a           (o_uart0_txd_a),
        .o_uart1_txdmasreq       (o_uart1_txdmasreq),
        .o_uart1_rxdmasreq       (o_uart1_rxdmasreq),
        .o_uart1_txdmabreq       (o_uart1_txdmabreq),
        .o_uart1_rxdmabreq       (o_uart1_rxdmabreq),
        .i_uart1_txdmaclr        (i_uart1_txdmaclr),
        .i_uart1_rxdmaclr        (i_uart1_rxdmaclr),
        .o_uart1_intr            (o_uart1_intr),
        .i_uart1_rxd_y           (i_uart1_rxd_y),
        .o_uart1_txd_a           (o_uart1_txd_a),
        .o_uart2_txdmasreq       (o_uart2_txdmasreq),
        .o_uart2_rxdmasreq       (o_uart2_rxdmasreq),
        .o_uart2_txdmabreq       (o_uart2_txdmabreq),
        .o_uart2_rxdmabreq       (o_uart2_rxdmabreq),
        .i_uart2_txdmaclr        (i_uart2_txdmaclr),
        .i_uart2_rxdmaclr        (i_uart2_rxdmaclr),
        .o_uart2_intr            (o_uart2_intr),
        .i_uart2_rxd_y           (i_uart2_rxd_y),
        .o_uart2_txd_a           (o_uart2_txd_a),
        .o_uart3_txdmasreq       (o_uart3_txdmasreq),
        .o_uart3_rxdmasreq       (o_uart3_rxdmasreq),
        .o_uart3_txdmabreq       (o_uart3_txdmabreq),
        .o_uart3_rxdmabreq       (o_uart3_rxdmabreq),
        .i_uart3_txdmaclr        (i_uart3_txdmaclr),
        .i_uart3_rxdmaclr        (i_uart3_rxdmaclr),
        .o_uart3_intr            (o_uart3_intr),
        .i_uart3_rxd_y           (i_uart3_rxd_y),
        .o_uart3_txd_a           (o_uart3_txd_a),
        .o_ssp0_intr             (o_ssp0_intr),
        .o_ssp0_txdamsreq        (o_ssp0_txdamsreq),
        .o_ssp0_rxdmasreq        (o_ssp0_rxdmasreq),
        .o_ssp0_txdmabreq        (o_ssp0_txdmabreq),
        .o_ssp0_rxdmabreq        (o_ssp0_rxdmabreq),
        .i_ssp0_txdmaclr         (i_ssp0_txdmaclr),
        .i_ssp0_rxdmaclr         (i_ssp0_rxdmaclr),
        .i_ssp0_clk_y            (i_ssp0_clk_y),
        .o_ssp0_clk_a            (o_ssp0_clk_a),
        .o_ssp0_clk_oe           (o_ssp0_clk_oe),
        .i_ssp0_csn_y            (i_ssp0_csn_y),
        .o_ssp0_csn_a            (o_ssp0_csn_a),
        .o_ssp0_csn_oe           (o_ssp0_csn_oe),
        .i_ssp0_rx_y             (i_ssp0_rx_y),
        .o_ssp0_tx_a             (o_ssp0_tx_a),
        .o_ssp1_intr             (o_ssp1_intr),
        .o_ssp1_txdamsreq        (o_ssp1_txdamsreq),
        .o_ssp1_rxdmasreq        (o_ssp1_rxdmasreq),
        .o_ssp1_txdmabreq        (o_ssp1_txdmabreq),
        .o_ssp1_rxdmabreq        (o_ssp1_rxdmabreq),
        .i_ssp1_txdmaclr         (i_ssp1_txdmaclr),
        .i_ssp1_rxdmaclr         (i_ssp1_rxdmaclr),
        .i_ssp1_clk_y            (i_ssp1_clk_y),
        .o_ssp1_clk_a            (o_ssp1_clk_a),
        .o_ssp1_clk_oe           (o_ssp1_clk_oe),
        .i_ssp1_csn_y            (i_ssp1_csn_y),
        .o_ssp1_csn_a            (o_ssp1_csn_a),
        .o_ssp1_csn_oe           (o_ssp1_csn_oe),
        .i_ssp1_rx_y             (i_ssp1_rx_y),
        .o_ssp1_tx_a             (o_ssp1_tx_a),
        .o_ssp2_intr             (o_ssp2_intr),
        .o_ssp2_txdamsreq        (o_ssp2_txdamsreq),
        .o_ssp2_rxdmasreq        (o_ssp2_rxdmasreq),
        .o_ssp2_txdmabreq        (o_ssp2_txdmabreq),
        .o_ssp2_rxdmabreq        (o_ssp2_rxdmabreq),
        .i_ssp2_txdmaclr         (i_ssp2_txdmaclr),
        .i_ssp2_rxdmaclr         (i_ssp2_rxdmaclr),
        .i_ssp2_clk_y            (i_ssp2_clk_y),
        .o_ssp2_clk_a            (o_ssp2_clk_a),
        .o_ssp2_clk_oe           (o_ssp2_clk_oe),
        .i_ssp2_csn_y            (i_ssp2_csn_y),
        .o_ssp2_csn_a            (o_ssp2_csn_a),
        .o_ssp2_csn_oe           (o_ssp2_csn_oe),
        .i_ssp2_rx_y             (i_ssp2_rx_y),
        .o_ssp2_tx_a             (o_ssp2_tx_a),
        .o_ssp3_intr             (o_ssp3_intr),
        .o_ssp3_txdamsreq        (o_ssp3_txdamsreq),
        .o_ssp3_rxdmasreq        (o_ssp3_rxdmasreq),
        .o_ssp3_txdmabreq        (o_ssp3_txdmabreq),
        .o_ssp3_rxdmabreq        (o_ssp3_rxdmabreq),
        .i_ssp3_txdmaclr         (i_ssp3_txdmaclr),
        .i_ssp3_rxdmaclr         (i_ssp3_rxdmaclr),
        .i_ssp3_clk_y            (i_ssp3_clk_y),
        .o_ssp3_clk_a            (o_ssp3_clk_a),
        .o_ssp3_clk_oe           (o_ssp3_clk_oe),
        .i_ssp3_csn_y            (i_ssp3_csn_y),
        .o_ssp3_csn_a            (o_ssp3_csn_a),
        .o_ssp3_csn_oe           (o_ssp3_csn_oe),
        .i_ssp3_rx_y             (i_ssp3_rx_y),
        .o_ssp3_tx_a             (o_ssp3_tx_a),
        .o_timer0_intr           (o_timer0_intr),
        .o_timer1_intr           (o_timer1_intr),
        .o_timer2_intr           (o_timer2_intr),
        .o_timer3_intr           (o_timer3_intr),
        .o_gpio0_intr            (o_gpio0_intr),
        .i_gpio0_y               (i_gpio0_y),
        .o_gpio0_a               (o_gpio0_a),
        .o_gpio0_oe              (o_gpio0_oe),
        .o_gpio1_intr            (o_gpio1_intr),
        .i_gpio1_y               (i_gpio1_y),
        .o_gpio1_a               (o_gpio1_a),
        .o_gpio1_oe              (o_gpio1_oe),
        .o_gpio2_intr            (o_gpio2_intr),
        .i_gpio2_y               (i_gpio2_y),
        .o_gpio2_a               (o_gpio2_a),
        .o_gpio2_oe              (o_gpio2_oe),
        .o_gpio3_intr            (o_gpio3_intr),
        .i_gpio3_y               (i_gpio3_y),
        .o_gpio3_a               (o_gpio3_a),
        .o_gpio3_oe              (o_gpio3_oe),
        .o_gpio4_intr            (o_gpio4_intr),
        .i_gpio4_y               (i_gpio4_y),
        .o_gpio4_a               (o_gpio4_a),
        .o_gpio4_oe              (o_gpio4_oe),
        .o_gpio5_intr            (o_gpio5_intr),
        .i_gpio5_y               (i_gpio5_y),
        .o_gpio5_a               (o_gpio5_a),
        .o_gpio5_oe              (o_gpio5_oe),
        .o_gpio6_intr            (o_gpio6_intr),
        .i_gpio6_y               (i_gpio6_y),
        .o_gpio6_a               (o_gpio6_a),
        .o_gpio6_oe              (o_gpio6_oe),
        .o_gpio7_intr            (o_gpio7_intr),
        .i_gpio7_y               (i_gpio7_y),
        .o_gpio7_a               (o_gpio7_a),
        .o_gpio7_oe              (o_gpio7_oe),
        .o_gpio8_intr            (o_gpio8_intr),
        .i_gpio8_y               (i_gpio8_y),
        .o_gpio8_a               (o_gpio8_a),
        .o_gpio8_oe              (o_gpio8_oe),
        .o_gpio9_intr            (o_gpio9_intr),
        .i_gpio9_y               (i_gpio9_y),
        .o_gpio9_a               (o_gpio9_a),
        .o_gpio9_oe              (o_gpio9_oe),
        .o_gpio10_intr           (o_gpio10_intr),
        .i_gpio10_y              (i_gpio10_y),
        .o_gpio10_a              (o_gpio10_a),
        .o_gpio10_oe             (o_gpio10_oe),
        .o_gpio11_intr           (o_gpio11_intr),
        .i_gpio11_y              (i_gpio11_y),
        .o_gpio11_a              (o_gpio11_a),
        .o_gpio11_oe             (o_gpio11_oe),
        .o_gpio12_intr           (o_gpio12_intr),
        .i_gpio12_y              (i_gpio12_y),
        .o_gpio12_a              (o_gpio12_a),
        .o_gpio12_oe             (o_gpio12_oe),
        .o_gpio13_intr           (o_gpio13_intr),
        .i_gpio13_y              (i_gpio13_y),
        .o_gpio13_a              (o_gpio13_a),
        .o_gpio13_oe             (o_gpio13_oe),
        .o_gpio14_intr           (o_gpio14_intr),
        .i_gpio14_y              (i_gpio14_y),
        .o_gpio14_a              (o_gpio14_a),
        .o_gpio14_oe             (o_gpio14_oe),
        .o_gpio15_intr           (o_gpio15_intr),
        .i_gpio15_y              (i_gpio15_y),
        .o_gpio15_a              (o_gpio15_a),
        .o_gpio15_oe             (o_gpio15_oe),
        .o_gpio16_intr           (o_gpio16_intr),
        .i_gpio16_y              (i_gpio16_y),
        .o_gpio16_a              (o_gpio16_a),
        .o_gpio16_oe             (o_gpio16_oe),
        .o_gpio17_intr           (o_gpio17_intr),
        .i_gpio17_y              (i_gpio17_y),
        .o_gpio17_a              (o_gpio17_a),
        .o_gpio17_oe             (o_gpio17_oe),
        .o_gpio18_intr           (o_gpio18_intr),
        .i_gpio18_y              (i_gpio18_y),
        .o_gpio18_a              (o_gpio18_a),
        .o_gpio18_oe             (o_gpio18_oe),
        .o_gpio19_intr           (o_gpio19_intr),
        .i_gpio19_y              (i_gpio19_y),
        .o_gpio19_a              (o_gpio19_a),
        .o_gpio19_oe             (o_gpio19_oe),
        .o_wdt_intr              (o_wdt_intr),
        .o_wdt_nresetout         (o_wdt_nresetout),
        .o_rtc_tic_irq0          (o_rtc_tic_irq0),
        .o_rtc_tic_irq1          (o_rtc_tic_irq1),
        .o_rtc_alarm_irq         (o_rtc_alarm_irq),
        .i_rtc_xin_ck            (i_rtc_xin_ck),
        .o_adc_clk               (o_adc_clk),
        .o_adc_pd                (o_adc_pd),
        .o_adc_soc               (o_adc_soc),
        .o_adc_sel               (o_adc_sel),
        .i_adc_eoc               (i_adc_eoc),
        .i_adc_data              (i_adc_data)
    );

    pnai70x_crm_peri u_crm_peri (
        .i_apb_pclk              (i_clk_peri_hpdf),
        .i_apb_prstn             (i_rstn_peri_hpdf),
        .i_apb_psel              (peri_sub_o_crm_apb_psel),
        .i_apb_penable           (peri_sub_o_crm_apb_penable),
        .i_apb_pwrite            (peri_sub_o_crm_apb_pwrite),
        .i_apb_paddr             (peri_sub_o_crm_apb_paddr),
        .i_apb_pwdata            (peri_sub_o_crm_apb_pwdata),
        .o_apb_prdata            (peri_sub_i_crm_apb_prdata),
        .i_rstn_peri_hpdf        (i_rstn_peri_hpdf),
        .i_clk_peri_hpdf         (i_clk_peri_hpdf),
        .i_clk_peri_codec        (i_clk_peri_codec),
        .i_i2s0_codck_y          (i_i2s0_codck_y),
        .i_i2s1_codck_y          (i_i2s1_codck_y),
        .o_clk_pclk_i2s0         (crm_peri_o_clk_pclk_i2s0),
        .o_rstn_pclk_i2s0        (crm_peri_o_rstn_pclk_i2s0),
        .o_clk_pclk_i2s1         (crm_peri_o_clk_pclk_i2s1),
        .o_rstn_pclk_i2s1        (crm_peri_o_rstn_pclk_i2s1),
        .o_clk_pclk_i2c0         (crm_peri_o_clk_pclk_i2c0),
        .o_rstn_pclk_i2c0        (crm_peri_o_rstn_pclk_i2c0),
        .o_clk_pclk_i2c1         (crm_peri_o_clk_pclk_i2c1),
        .o_rstn_pclk_i2c1        (crm_peri_o_rstn_pclk_i2c1),
        .o_clk_pclk_i2c2         (crm_peri_o_clk_pclk_i2c2),
        .o_rstn_pclk_i2c2        (crm_peri_o_rstn_pclk_i2c2),
        .o_clk_pclk_i2c3         (crm_peri_o_clk_pclk_i2c3),
        .o_rstn_pclk_i2c3        (crm_peri_o_rstn_pclk_i2c3),
        .o_clk_pclk_uart0        (crm_peri_o_clk_pclk_uart0),
        .o_rstn_pclk_uart0       (crm_peri_o_rstn_pclk_uart0),
        .o_clk_pclk_uart1        (crm_peri_o_clk_pclk_uart1),
        .o_rstn_pclk_uart1       (crm_peri_o_rstn_pclk_uart1),
        .o_clk_pclk_uart2        (crm_peri_o_clk_pclk_uart2),
        .o_rstn_pclk_uart2       (crm_peri_o_rstn_pclk_uart2),
        .o_clk_pclk_uart3        (crm_peri_o_clk_pclk_uart3),
        .o_rstn_pclk_uart3       (crm_peri_o_rstn_pclk_uart3),
        .o_clk_pclk_spi0         (crm_peri_o_clk_pclk_spi0),
        .o_rstn_pclk_spi0        (crm_peri_o_rstn_pclk_spi0),
        .o_clk_pclk_spi1         (crm_peri_o_clk_pclk_spi1),
        .o_rstn_pclk_spi1        (crm_peri_o_rstn_pclk_spi1),
        .o_clk_pclk_spi2         (crm_peri_o_clk_pclk_spi2),
        .o_rstn_pclk_spi2        (crm_peri_o_rstn_pclk_spi2),
        .o_clk_pclk_spi3         (crm_peri_o_clk_pclk_spi3),
        .o_rstn_pclk_spi3        (crm_peri_o_rstn_pclk_spi3),
        .o_clk_pclk_timer0       (crm_peri_o_clk_pclk_timer0),
        .o_rstn_pclk_timer0      (crm_peri_o_rstn_pclk_timer0),
        .o_clk_pclk_timer1       (crm_peri_o_clk_pclk_timer1),
        .o_rstn_pclk_timer1      (crm_peri_o_rstn_pclk_timer1),
        .o_clk_pclk_timer2       (crm_peri_o_clk_pclk_timer2),
        .o_rstn_pclk_timer2      (crm_peri_o_rstn_pclk_timer2),
        .o_clk_pclk_timer3       (crm_peri_o_clk_pclk_timer3),
        .o_rstn_pclk_timer3      (crm_peri_o_rstn_pclk_timer3),
        .o_clk_pclk_gpio0        (crm_peri_o_clk_pclk_gpio0),
        .o_rstn_pclk_gpio0       (crm_peri_o_rstn_pclk_gpio0),
        .o_clk_pclk_gpio1        (crm_peri_o_clk_pclk_gpio1),
        .o_rstn_pclk_gpio1       (crm_peri_o_rstn_pclk_gpio1),
        .o_clk_pclk_gpio2        (crm_peri_o_clk_pclk_gpio2),
        .o_rstn_pclk_gpio2       (crm_peri_o_rstn_pclk_gpio2),
        .o_clk_pclk_gpio3        (crm_peri_o_clk_pclk_gpio3),
        .o_rstn_pclk_gpio3       (crm_peri_o_rstn_pclk_gpio3),
        .o_clk_pclk_gpio4        (crm_peri_o_clk_pclk_gpio4),
        .o_rstn_pclk_gpio4       (crm_peri_o_rstn_pclk_gpio4),
        .o_clk_pclk_gpio5        (crm_peri_o_clk_pclk_gpio5),
        .o_rstn_pclk_gpio5       (crm_peri_o_rstn_pclk_gpio5),
        .o_clk_pclk_gpio6        (crm_peri_o_clk_pclk_gpio6),
        .o_rstn_pclk_gpio6       (crm_peri_o_rstn_pclk_gpio6),
        .o_clk_pclk_gpio7        (crm_peri_o_clk_pclk_gpio7),
        .o_rstn_pclk_gpio7       (crm_peri_o_rstn_pclk_gpio7),
        .o_clk_pclk_gpio8        (crm_peri_o_clk_pclk_gpio8),
        .o_rstn_pclk_gpio8       (crm_peri_o_rstn_pclk_gpio8),
        .o_clk_pclk_gpio9        (crm_peri_o_clk_pclk_gpio9),
        .o_rstn_pclk_gpio9       (crm_peri_o_rstn_pclk_gpio9),
        .o_clk_pclk_gpio10       (crm_peri_o_clk_pclk_gpio10),
        .o_rstn_pclk_gpio10      (crm_peri_o_rstn_pclk_gpio10),
        .o_clk_pclk_gpio11       (crm_peri_o_clk_pclk_gpio11),
        .o_rstn_pclk_gpio11      (crm_peri_o_rstn_pclk_gpio11),
        .o_clk_pclk_gpio12       (crm_peri_o_clk_pclk_gpio12),
        .o_rstn_pclk_gpio12      (crm_peri_o_rstn_pclk_gpio12),
        .o_clk_pclk_gpio13       (crm_peri_o_clk_pclk_gpio13),
        .o_rstn_pclk_gpio13      (crm_peri_o_rstn_pclk_gpio13),
        .o_clk_pclk_gpio14       (crm_peri_o_clk_pclk_gpio14),
        .o_rstn_pclk_gpio14      (crm_peri_o_rstn_pclk_gpio14),
        .o_clk_pclk_gpio15       (crm_peri_o_clk_pclk_gpio15),
        .o_rstn_pclk_gpio15      (crm_peri_o_rstn_pclk_gpio15),
        .o_clk_pclk_gpio16       (crm_peri_o_clk_pclk_gpio16),
        .o_rstn_pclk_gpio16      (crm_peri_o_rstn_pclk_gpio16),
        .o_clk_pclk_gpio17       (crm_peri_o_clk_pclk_gpio17),
        .o_rstn_pclk_gpio17      (crm_peri_o_rstn_pclk_gpio17),
        .o_clk_pclk_gpio18       (crm_peri_o_clk_pclk_gpio18),
        .o_rstn_pclk_gpio18      (crm_peri_o_rstn_pclk_gpio18),
        .o_clk_pclk_gpio19       (crm_peri_o_clk_pclk_gpio19),
        .o_rstn_pclk_gpio19      (crm_peri_o_rstn_pclk_gpio19),
        .o_clk_pclk_wdt          (crm_peri_o_clk_pclk_wdt),
        .o_rstn_pclk_wdt         (crm_peri_o_rstn_pclk_wdt),
        .o_clk_pclk_rtc          (crm_peri_o_clk_pclk_rtc),
        .o_rstn_pclk_rtc         (crm_peri_o_rstn_pclk_rtc),
        .o_clk_pclk_adc          (crm_peri_o_clk_pclk_adc),
        .o_rstn_pclk_adc         (crm_peri_o_rstn_pclk_adc),
        .o_clk_peri_bus          (crm_peri_o_clk_peri_bus),
        .o_rstn_peri_bus         (crm_peri_o_rstn_peri_bus),
        .o_clk_codec_clk0        (crm_peri_o_clk_codec_clk0),
        .o_clk_codec_clk1        (crm_peri_o_clk_codec_clk1),
        .i_scan_clk              (i_test_clk),
        .i_scan_mode             (i_test_mode),
        .i_scan_rstn             (1'h0)
    );

endmodule