module bus_top (
    input           bclk   ,
    input           bresetn,
    // SI0
    input           s0_psel    ,
    input           s0_penable ,
    input  [31:0]   s0_paddr   ,
    input           s0_pwrite  ,
    input  [31:0]   s0_pwdata  ,
    input  [2:0]    s0_pprot   ,
    input  [3:0]    s0_pstrb   ,
    output [31:0]   s0_prdata  ,
    output          s0_pready  ,
    output          s0_pslverr ,
    // SI1
    input  [1:0]     s1_htrans   ,
    input  [31:0    s1_haddr    ,
    input           s1_hwrite   ,
    input  [2:0]    s1_hsize    ,
    input  [2:0]    s1_hburst   ,
    input  [1:0]    s1_hwdata   ,
    input           s1_hmastlock,
    output [31:0]   s1_hrdata   ,
    output          s1_hready   ,
    output [1:0]    s1_hresp    ,
    // SI2
    input  [3:0]    s2_awid     ,
    input  [31:0]   s2_awaddr   ,
    input  [3:0]    s2_awlen    ,
    input  [2:0]    s2_awsize   ,
    input  [1:0]    s2_awburst  ,
    input  [1:0]    s2_awlock   ,
    input  [3:0]    s2_awcache  ,
    input  [2:0]    s2_awprot   ,
    input           s2_awvalid  ,
    output          s2_awready  ,
    input  [3:0]    s2_wid      ,
    input  [127:0]  s2_wdata    ,
    input  [15:0]   s2_wstrb    ,
    input           s2_wlast    ,
    input           s2_wvalid   ,
    output          s2_wready   ,
    output [3:0]    s2_bid      ,
    output [1:0]    s2_bresp    ,
    output          s2_bvalid   ,
    input           s2_bready   ,
    input  [3:0]    s2_arid     ,
    input  [31:0]   s2_araddr   ,
    input  [3:0]    s2_arlen    ,
    input  [2:0]    s2_arsize   ,
    input  [1:0]    s2_arburst  ,
    input  [1:0]    s2_arlock   ,
    input  [3:0]    s2_arcache  ,
    input  [2:0]    s2_arprot   ,
    input           s2_arvalid  ,
    output          s2_arready  ,
    output [3:0]    s2_rid      ,
    output [127:0]  s2_rdata    ,
    output [1:0]    s2_rresp    ,
    output          s2_rlast    ,
    output          s2_rvalid   ,
    input           s2_rready   ,
    // MI0 - 
    output          mi0_psel    ,
    output          mi0_penable ,
    output [31:0]   mi0_paddr   ,
    output          mi0_pwrite  ,
    output [31:0]   mi0_pwdata  ,
    output [2:0]    mi0_pprot   ,
    output [3:0]    mi0_pstrb   ,
    input  [31:0]   mi0_prdata  ,
    input           mi0_pready  ,
    input           mi0_pslverr ,
    // MI1
    output [1:0     mi1_htrans   ,
    output [31:0    mi1_haddr    ,
    output          mi1_hwrite   ,
    output [2:0]    mi1_hsize    ,
    output [2:0]    mi1_hburst   ,
    output [1:0]    mi1_hwdata   ,
    output          mi1_hmastlock,
    input  [31:0]   mi1_hrdata   ,
    input           mi1_hready   ,
    input  [1:0]    mi1_hresp    ,
    // MI2
    output [3:0]    mi2_awid   ,
    output [31:0]   mi2_awaddr ,
    output [3:0]    mi2_awlen  ,
    output [2:0]    mi2_awsize ,
    output [1:0]    mi2_awburst,
    output [1:0]    mi2_awlock ,
    output [3:0]    mi2_awcache,
    output [2:0]    mi2_awprot ,
    output          mi2_awvalid,
    input           mi2_awready,
    output [3:0]    mi2_wid    ,
    output [127:0]  mi2_wdata  ,
    output [15:0]   mi2_wstrb  ,
    output          mi2_wlast  ,
    output          mi2_wvalid ,
    input           mi2_wready ,
    input  [3:0]    mi2_bid    ,
    input  [1:0]    mi2_bresp  ,
    input           mi2_bvalid ,
    output          mi2_bready ,
    output [3:0]    mi2_arid   ,
    output [31:0]   mi2_araddr ,
    output [3:0]    mi2_arlen  ,
    output [2:0]    mi2_arsize ,
    output [1:0]    mi2_arburst,
    output [1:0]    mi2_arlock ,
    output [3:0]    mi2_arcache,
    output [2:0]    mi2_arprot ,
    output          mi2_arvalid,
    input           mi2_arready,
    input  [3:0]    mi2_rid    ,
    input  [127:0]  mi2_rdata  ,
    input  [1:0]    mi2_rresp  ,
    input           mi2_rlast  ,
    input           mi2_rvalid ,
    output          mi2_rready 
);

endmodule