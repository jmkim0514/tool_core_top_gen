//==============================================================================
//
// Project : MVP
//
// Verilog RTL(Behavioral) model
//
// This confidential and proprietary source code may be used only as authorized
// by a licensing agreement from ALPHAHOLDINGS Limited. The entire notice above
// must be reproduced on all authorized copies and copies may only be made to
// the extent permitted by a licensing agreement from ALPHAHOLDINGS Limited.
//
// COPYRIGHT (C) ALPHAHOLDINGS, inc. 2022
//
//==============================================================================
// File name : keti_hpdf
// Version : v1.1
// Description :
// Simulator : NC Verilog
// Created by : syhan
// Date : 2023-09-21  17:31
//==============================================================================

module keti_hpdf (
    input              i_test_bypass,
    input              i_rstn_peri2keti,
    input              i_clk_peri2keti,
    input              i_clk_keti_ip,
    input              i_scan_clk,
    input              i_scan_mode,
    input              i_test_rstn,
    input              i_test_mode,
    output             o_irq_keti,
    input   [ 38:  0]  i_ema,
    input   [ 31:  0]  i_paddr_peri2keti_m3,
    input              i_pwrite_peri2keti_m3,
    input              i_pselx_peri2keti_m3,
    input              i_penable_peri2keti_m3,
    input   [ 31:  0]  i_pwdata_peri2keti_m3,
    output             o_pready_peri2keti_m3,
    output  [ 31:  0]  o_prdata_peri2keti_m3,
    output             o_pslverr_peri2keti_m3,
    output  [  1:  0]  o_arid_keti2main_0,
    output  [  7:  0]  o_arlen_keti2main_0,
    output  [  2:  0]  o_arsize_keti2main_0,
    output  [  1:  0]  o_arburst_keti2main_0,
    output             o_arlock_keti2main_0,
    output  [  3:  0]  o_arcache_keti2main_0,
    output  [  2:  0]  o_arprot_keti2main_0,
    output  [ 31:  0]  o_araddr_keti2main_0,
    output             o_arvalid_keti2main_0,
    input              i_arready_keti2main_0,
    input   [  1:  0]  i_rid_keti2main_0,
    input              i_rvalid_keti2main_0,
    input   [ 63:  0]  i_rdata_keti2main_0,
    input              i_rlast_keti2main_0,
    output             o_rready_keti2main_0,
    input   [  1:  0]  i_rresp_keti2main_0,
    output  [  1:  0]  o_awid_keti2main_0,
    output  [  7:  0]  o_awlen_keti2main_0,
    output  [  2:  0]  o_awsize_keti2main_0,
    output  [  1:  0]  o_awburst_keti2main_0,
    output             o_awlock_keti2main_0,
    output  [  3:  0]  o_awcache_keti2main_0,
    output  [  2:  0]  o_awprot_keti2main_0,
    output  [ 31:  0]  o_awaddr_keti2main_0,
    output             o_awvalid_keti2main_0,
    input              i_awready_keti2main_0,
    output  [ 63:  0]  o_wdata_keti2main_0,
    output  [  7:  0]  o_wstrb_keti2main_0,
    output             o_wlast_keti2main_0,
    output             o_wvalid_keti2main_0,
    input              i_wready_keti2main_0,
    input   [  1:  0]  i_bresp_keti2main_0,
    input   [  1:  0]  i_bid_keti2main_0,
    input              i_bvalid_keti2main_0,
    output             o_bready_keti2main_0,
    output  [  1:  0]  o_awuser_keti2main_0,
    output  [  1:  0]  o_aruser_keti2main_0,
    output  [  2:  0]  o_arid_keti2main_1,
    output  [  7:  0]  o_arlen_keti2main_1,
    output  [  2:  0]  o_arsize_keti2main_1,
    output  [  1:  0]  o_arburst_keti2main_1,
    output             o_arlock_keti2main_1,
    output  [  3:  0]  o_arcache_keti2main_1,
    output  [  2:  0]  o_arprot_keti2main_1,
    output  [ 31:  0]  o_araddr_keti2main_1,
    output             o_arvalid_keti2main_1,
    input              i_arready_keti2main_1,
    input   [  2:  0]  i_rid_keti2main_1,
    input              i_rvalid_keti2main_1,
    input   [127:  0]  i_rdata_keti2main_1,
    input              i_rlast_keti2main_1,
    output             o_rready_keti2main_1,
    input   [  1:  0]  i_rresp_keti2main_1,
    output  [  2:  0]  o_awid_keti2main_1,
    output  [  7:  0]  o_awlen_keti2main_1,
    output  [  2:  0]  o_awsize_keti2main_1,
    output  [  1:  0]  o_awburst_keti2main_1,
    output             o_awlock_keti2main_1,
    output  [  3:  0]  o_awcache_keti2main_1,
    output  [  2:  0]  o_awprot_keti2main_1,
    output  [ 31:  0]  o_awaddr_keti2main_1,
    output             o_awvalid_keti2main_1,
    input              i_awready_keti2main_1,
    output  [127:  0]  o_wdata_keti2main_1,
    output  [ 15:  0]  o_wstrb_keti2main_1,
    output             o_wlast_keti2main_1,
    output             o_wvalid_keti2main_1,
    input              i_wready_keti2main_1,
    input   [  2:  0]  i_bid_keti2main_1,
    input   [  1:  0]  i_bresp_keti2main_1,
    input              i_bvalid_keti2main_1,
    output             o_bready_keti2main_1,
    output  [  1:  0]  o_awuser_keti2main_1,
    output  [  1:  0]  o_aruser_keti2main_1
);

    wire            keti_crm_o_clk_keti_peri;
    wire            keti_crm_o_rstn_keti_peri;
    wire            keti_crm_o_clk_keti_ip;
    wire            keti_crm_o_rstn_keti_ip;
    wire            keti_sub_o_psel_keti_crm;
    wire            keti_sub_o_penable_keti_crm;
    wire            keti_sub_o_pwrite_keti_crm;
    wire    [11:0]  keti_sub_o_paddr_keti_crm;
    wire    [31:0]  keti_sub_o_pwdata_keti_crm;
    wire    [31:0]  keti_sub_i_prdata_keti_crm;


    mvp_crm_keti u_keti_crm (
        .i_test_bypass            (i_test_bypass),
        .i_rstn_keti_crm          (i_rstn_peri2keti),
        .i_apb_pclk               (i_clk_peri2keti),
        .i_apb_prstn              (i_rstn_peri2keti),
        .i_apb_psel               (keti_sub_o_psel_keti_crm),
        .i_apb_penable            (keti_sub_o_penable_keti_crm),
        .i_apb_pwrite             (keti_sub_o_pwrite_keti_crm),
        .i_apb_paddr              (keti_sub_o_paddr_keti_crm),
        .i_apb_pwdata             (keti_sub_o_pwdata_keti_crm),
        .o_apb_prdata             (keti_sub_i_prdata_keti_crm),
        .i_clk_peri2keti          (i_clk_peri2keti),
        .i_clk_keti_ip            (i_clk_keti_ip),
        .o_clk_keti_peri          (keti_crm_o_clk_keti_peri),
        .o_rstn_keti_peri         (keti_crm_o_rstn_keti_peri),
        .o_clk_keti_ip            (keti_crm_o_clk_keti_ip),
        .o_rstn_keti_ip           (keti_crm_o_rstn_keti_ip),
        .i_scan_clk               (i_scan_clk),
        .i_scan_mode              (i_scan_mode),
        .i_scan_rstn              (i_test_rstn)
    );

    keti_sub u_keti_sub (
        .i_clk_keti_peri          (keti_crm_o_clk_keti_peri),
        .i_rstn_keti_peri         (keti_crm_o_rstn_keti_peri),
        .i_clk_keti_sfr           (keti_crm_o_clk_keti_ip),
        .i_rstn_keti_sfr          (keti_crm_o_rstn_keti_ip),
        .i_clk_keti_ip            (keti_crm_o_clk_keti_ip),
        .i_rstn_keti_ip           (keti_crm_o_rstn_keti_ip),
        .i_paddr_peri2keti_m3     (i_paddr_peri2keti_m3),
        .i_pwrite_peri2keti_m3    (i_pwrite_peri2keti_m3),
        .i_pselx_peri2keti_m3     (i_pselx_peri2keti_m3),
        .i_penable_peri2keti_m3   (i_penable_peri2keti_m3),
        .i_pwdata_peri2keti_m3    (i_pwdata_peri2keti_m3),
        .o_pready_peri2keti_m3    (o_pready_peri2keti_m3),
        .o_prdata_peri2keti_m3    (o_prdata_peri2keti_m3),
        .o_pslverr_peri2keti_m3   (o_pslverr_peri2keti_m3),
        .o_psel_keti_crm          (keti_sub_o_psel_keti_crm),
        .o_penable_keti_crm       (keti_sub_o_penable_keti_crm),
        .o_pwrite_keti_crm        (keti_sub_o_pwrite_keti_crm),
        .o_paddr_keti_crm         (keti_sub_o_paddr_keti_crm),
        .o_pwdata_keti_crm        (keti_sub_o_pwdata_keti_crm),
        .i_prdata_keti_crm        (keti_sub_i_prdata_keti_crm),
        .o_arid_keti2main_0       (o_arid_keti2main_0),
        .o_arlen_keti2main_0      (o_arlen_keti2main_0),
        .o_arsize_keti2main_0     (o_arsize_keti2main_0),
        .o_arburst_keti2main_0    (o_arburst_keti2main_0),
        .o_arlock_keti2main_0     (o_arlock_keti2main_0),
        .o_arcache_keti2main_0    (o_arcache_keti2main_0),
        .o_arprot_keti2main_0     (o_arprot_keti2main_0),
        .o_araddr_keti2main_0     (o_araddr_keti2main_0),
        .o_arvalid_keti2main_0    (o_arvalid_keti2main_0),
        .i_arready_keti2main_0    (i_arready_keti2main_0),
        .i_rid_keti2main_0        (i_rid_keti2main_0),
        .i_rvalid_keti2main_0     (i_rvalid_keti2main_0),
        .i_rdata_keti2main_0      (i_rdata_keti2main_0),
        .i_rlast_keti2main_0      (i_rlast_keti2main_0),
        .o_rready_keti2main_0     (o_rready_keti2main_0),
        .i_rresp_keti2main_0      (i_rresp_keti2main_0),
        .o_awid_keti2main_0       (o_awid_keti2main_0),
        .o_awlen_keti2main_0      (o_awlen_keti2main_0),
        .o_awsize_keti2main_0     (o_awsize_keti2main_0),
        .o_awburst_keti2main_0    (o_awburst_keti2main_0),
        .o_awlock_keti2main_0     (o_awlock_keti2main_0),
        .o_awcache_keti2main_0    (o_awcache_keti2main_0),
        .o_awprot_keti2main_0     (o_awprot_keti2main_0),
        .o_awaddr_keti2main_0     (o_awaddr_keti2main_0),
        .o_awvalid_keti2main_0    (o_awvalid_keti2main_0),
        .i_awready_keti2main_0    (i_awready_keti2main_0),
        .o_wdata_keti2main_0      (o_wdata_keti2main_0),
        .o_wstrb_keti2main_0      (o_wstrb_keti2main_0),
        .o_wlast_keti2main_0      (o_wlast_keti2main_0),
        .o_wvalid_keti2main_0     (o_wvalid_keti2main_0),
        .i_wready_keti2main_0     (i_wready_keti2main_0),
        .i_bresp_keti2main_0      (i_bresp_keti2main_0),
        .i_bid_keti2main_0        (i_bid_keti2main_0),
        .i_bvalid_keti2main_0     (i_bvalid_keti2main_0),
        .o_bready_keti2main_0     (o_bready_keti2main_0),
        .o_awuser_keti2main_0     (o_awuser_keti2main_0),
        .o_aruser_keti2main_0     (o_aruser_keti2main_0),
        .o_arid_keti2main_1       (o_arid_keti2main_1),
        .o_arlen_keti2main_1      (o_arlen_keti2main_1),
        .o_arsize_keti2main_1     (o_arsize_keti2main_1),
        .o_arburst_keti2main_1    (o_arburst_keti2main_1),
        .o_arlock_keti2main_1     (o_arlock_keti2main_1),
        .o_arcache_keti2main_1    (o_arcache_keti2main_1),
        .o_arprot_keti2main_1     (o_arprot_keti2main_1),
        .o_araddr_keti2main_1     (o_araddr_keti2main_1),
        .o_arvalid_keti2main_1    (o_arvalid_keti2main_1),
        .i_arready_keti2main_1    (i_arready_keti2main_1),
        .i_rid_keti2main_1        (i_rid_keti2main_1),
        .i_rvalid_keti2main_1     (i_rvalid_keti2main_1),
        .i_rdata_keti2main_1      (i_rdata_keti2main_1),
        .i_rlast_keti2main_1      (i_rlast_keti2main_1),
        .o_rready_keti2main_1     (o_rready_keti2main_1),
        .i_rresp_keti2main_1      (i_rresp_keti2main_1),
        .o_awid_keti2main_1       (o_awid_keti2main_1),
        .o_awlen_keti2main_1      (o_awlen_keti2main_1),
        .o_awsize_keti2main_1     (o_awsize_keti2main_1),
        .o_awburst_keti2main_1    (o_awburst_keti2main_1),
        .o_awlock_keti2main_1     (o_awlock_keti2main_1),
        .o_awcache_keti2main_1    (o_awcache_keti2main_1),
        .o_awprot_keti2main_1     (o_awprot_keti2main_1),
        .o_awaddr_keti2main_1     (o_awaddr_keti2main_1),
        .o_awvalid_keti2main_1    (o_awvalid_keti2main_1),
        .i_awready_keti2main_1    (i_awready_keti2main_1),
        .o_wdata_keti2main_1      (o_wdata_keti2main_1),
        .o_wstrb_keti2main_1      (o_wstrb_keti2main_1),
        .o_wlast_keti2main_1      (o_wlast_keti2main_1),
        .o_wvalid_keti2main_1     (o_wvalid_keti2main_1),
        .i_wready_keti2main_1     (i_wready_keti2main_1),
        .i_bid_keti2main_1        (i_bid_keti2main_1),
        .i_bresp_keti2main_1      (i_bresp_keti2main_1),
        .i_bvalid_keti2main_1     (i_bvalid_keti2main_1),
        .o_bready_keti2main_1     (o_bready_keti2main_1),
        .o_awuser_keti2main_1     (o_awuser_keti2main_1),
        .o_aruser_keti2main_1     (o_aruser_keti2main_1),
        .i_keti_test_mode         (i_test_mode),
        .o_irq_keti               (o_irq_keti),
        .i_ema                    (i_ema)
    );

endmodule